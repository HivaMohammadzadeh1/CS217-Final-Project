
//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 02:51:36 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [168:0] this_dat;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [127:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_dat[127:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_dat[151:128];
  wire  nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_dat[168];
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd128)) data_data_rsci (
      .d(nl_data_data_rsci_d[127:0]),
      .z(data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d),
      .z(data_rw_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd154),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [168:0] this_dat;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 02:51:31 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [137:0] this_dat;
  output [127:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [127:0] nl_data_data_data_rsci_d;
  assign nl_data_data_data_rsci_d = this_dat[127:0];
  wire [7:0] nl_data_logical_addr_rsci_d;
  assign nl_data_logical_addr_rsci_d = this_dat[137:130];
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd7),
  .width(32'sd128)) data_data_data_rsci (
      .d(nl_data_data_data_rsci_d[127:0]),
      .z(data_data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd9),
  .width(32'sd8)) data_logical_addr_rsci (
      .d(nl_data_logical_addr_rsci_d[7:0]),
      .z(data_logical_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd11),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd153),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [137:0] this_dat;
  output [127:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_data_rsc_z(data_data_data_rsc_z),
      .data_logical_addr_rsc_z(data_logical_addr_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 02:51:28 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [255:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [16:0] m_data_buf_240_0_lpi_1_dfm_240_224;
  reg [16:0] m_data_buf_240_0_lpi_1_dfm_208_192;
  reg [16:0] m_data_buf_240_0_lpi_1_dfm_176_160;
  reg [16:0] m_data_buf_240_0_lpi_1_dfm_144_128;
  reg [16:0] m_data_buf_240_0_lpi_1_dfm_112_96;
  reg [16:0] m_data_buf_240_0_lpi_1_dfm_80_64;
  reg [16:0] m_data_buf_240_0_lpi_1_dfm_48_32;
  reg [16:0] m_data_buf_240_0_lpi_1_dfm_16_0;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd13),
  .width(32'sd256)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd152),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd156)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = {15'b000000000000000 , m_data_buf_240_0_lpi_1_dfm_240_224 , 15'b000000000000000
      , m_data_buf_240_0_lpi_1_dfm_208_192 , 15'b000000000000000 , m_data_buf_240_0_lpi_1_dfm_176_160
      , 15'b000000000000000 , m_data_buf_240_0_lpi_1_dfm_144_128 , 15'b000000000000000
      , m_data_buf_240_0_lpi_1_dfm_112_96 , 15'b000000000000000 , m_data_buf_240_0_lpi_1_dfm_80_64
      , 15'b000000000000000 , m_data_buf_240_0_lpi_1_dfm_48_32 , 15'b000000000000000
      , m_data_buf_240_0_lpi_1_dfm_16_0};
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_240_0_lpi_1_dfm_240_224 <= 17'b00000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_240_0_lpi_1_dfm_240_224 <= m_data_rsci_idat[240:224];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_240_0_lpi_1_dfm_208_192 <= 17'b00000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_240_0_lpi_1_dfm_208_192 <= m_data_rsci_idat[208:192];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_240_0_lpi_1_dfm_176_160 <= 17'b00000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_240_0_lpi_1_dfm_176_160 <= m_data_rsci_idat[176:160];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_240_0_lpi_1_dfm_144_128 <= 17'b00000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_240_0_lpi_1_dfm_144_128 <= m_data_rsci_idat[144:128];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_240_0_lpi_1_dfm_112_96 <= 17'b00000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_240_0_lpi_1_dfm_112_96 <= m_data_rsci_idat[112:96];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_240_0_lpi_1_dfm_80_64 <= 17'b00000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_240_0_lpi_1_dfm_80_64 <= m_data_rsci_idat[80:64];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_240_0_lpi_1_dfm_48_32 <= 17'b00000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_240_0_lpi_1_dfm_48_32 <= m_data_rsci_idat[48:32];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_240_0_lpi_1_dfm_16_0 <= 17'b00000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_240_0_lpi_1_dfm_16_0 <= m_data_rsci_idat[16:0];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 01:32:50 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd15),
  .width(32'sd1)) data_rsci (
      .d(this_dat),
      .z(data_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd17),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd151),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 02:51:33 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [127:0] this_dat;
  reg [127:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [127:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd18),
  .width(32'sd128)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd150),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd155)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [127:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_mgc_muladd1_beh.v 
//muladd1
module PECore_mgc_muladd1(a,b,c,cst,d,z);
  // operation is z = a * (b + d) + c + cst
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_cst = 0;
  parameter signd_cst = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_axb = 1;
  parameter add_c = 1;
  parameter add_d = 1;
  parameter use_const = 1;

  function integer is_square_op;
    input integer alen;
  begin
    if (alen > 1) is_square_op = 0;
    else       is_square_op = 1;
  end endfunction

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_cst-1:0] cst; // spyglass disable SYNTH_5121,W240
  input  [width_d-1:0] d;
  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa;
  reg [width_b-signd_b:0] bb;
  reg [width_c-signd_c:0] cc;
  reg [width_d-signd_d:0] dd;
  reg [width_cst-signd_cst:0] cstin;

  localparam width_bd = (width_d) ? 1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b
                                                                          : width_d - signd_d)
                                  : width_b - signd_b;
  localparam is_square = is_square_op(width_a);
  localparam axb_len = (is_square)?width_bd+1+width_bd+1:width_a-signd_a+1+width_bd+1;

  reg [width_bd:0] bd;
  reg [axb_len-1:0] axb;



  // make all inputs signed
  always @(*) aa = signd_a ? a : {1'b0, a};
  always @(*) bb = signd_b ? b : {1'b0, b};
  generate if (width_c != 0) begin
    always @(*) cc = signd_c ? c : {1'b0, c};
  end endgenerate

  generate if (width_d) begin
    if ( !is_square) begin
      (* keep ="true" *) reg [width_d-signd_d:0] d_keep;
      always @(*) d_keep = signd_d ? d : {1'b0, d};
      always @(*) dd = d_keep;
    end else begin
      always @(*) dd = signd_d ? d : {1'b0, d};
    end
  end endgenerate

  always @(*) cstin = signd_cst ? cst : {1'b0, cst};

  // perform pre-adder
  generate
    if (width_d != 0) begin
      if (add_d) begin always @(*)  bd = $signed(bb) + $signed(dd); end
      else       begin always @(*)  bd = $signed(bb) - $signed(dd); end
    end else     begin always @(*)  bd = $signed(bb); end
  endgenerate

  generate
    if (is_square)
      always @(*) axb = $signed(bd) * $signed(bd);
    else
      always @(*) axb = $signed(aa) * $signed(bd);
  endgenerate

  // perform muladd1
  wire [width_z-1:0]  zz;

  generate
    if (use_const) begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc) + $signed(cstin); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc) + $signed(cstin); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb) + $signed(cstin); end else
      if (!add_axb && !add_c && width_c) begin assign zz = $signed(cstin) - $signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb) + $signed(cstin); end else
                                         begin assign zz = $signed(cstin) - $signed(axb); end
    end  else begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb); end else
      if (!add_axb && !add_c && width_c) begin assign zz = -$signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb); end else
                                         begin assign zz = -$signed(axb); end
    end
  endgenerate

  // adjust output
  assign z = zz;
endmodule // mgc_muladd1

//------> ./PECore_mgc_shift_l_beh_v5.v 
module PECore_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./PECore_mgc_mul2add1_pipe_beh.v 
//muladd1
module PECore_mgc_mul2add1_pipe(a,b,b2,c,d,d2,cst,clk,en,a_rst,s_rst,z);
  parameter gentype = 0;
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_b2 = 0;
  parameter signd_b2 = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_d2 = 0;
  parameter signd_d2 = 0;
  parameter width_e = 0;
  parameter signd_e = 0;
  parameter width_z = 0;
  parameter isadd = 1;
  parameter add_b2 = 1;
  parameter add_d2 = 1;
  parameter use_const = 1;
  parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
  parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
  parameter    a_rst_active =  1'b1;  // unused
  parameter    s_rst_active =  1'b1;  // unused
  parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
  parameter integer n_inreg = 32'd0;  // number of input registers

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_b2-1:0] b2; // spyglass disable SYNTH_5121,W240
  input  [width_c-1:0] c;
  input  [width_d-1:0] d;
  input  [width_d2-1:0] d2; // spyglass disable SYNTH_5121,W240
  input  [width_e-1:0] cst; // spyglass disable SYNTH_5121,W240

  input                clk;    // clock
  input                en;     // enable
  input                a_rst;  // spyglass disable SYNTH_5121,W240
  input                s_rst;  // spyglass disable SYNTH_5121,W240

  output [width_z-1:0] z;

  function integer MIN;
    input integer a, b;
  begin
    if (a > b) MIN = b;
    else       MIN = a;
  end endfunction

  function integer f_axb_stages;
    input integer gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d;
  begin
    if (gentype%2==0) begin
      if ((n_inreg > 1) && (width_a>18 | width_b>=19+signd_b | width_c>18 | width_d>=19+signd_d ))
        f_axb_stages = 1;
      else
        f_axb_stages = 0;
    end else begin
      if (n_inreg>1)
        f_axb_stages = 1;
      else
        f_axb_stages = 0;
    end
  end endfunction

  function integer f_cxd_stages;
    input integer gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d;
  begin
    if (gentype%2==0) begin
      f_cxd_stages = 0;
    end else begin
      if (n_inreg>1)
        f_cxd_stages = MIN(n_inreg-1,3);
      else
        f_cxd_stages = 0;
    end
  end endfunction

  function integer f_preadd_stages;
    input integer gentype,n_inreg,width_preaddin;
  begin
    if (gentype%2==0) begin
      f_preadd_stages = 0;
    end else begin
      if (n_inreg>1) begin
        if (width_preaddin>0)
          f_preadd_stages = 1;
        else
          f_preadd_stages = 0;
      end else
        f_preadd_stages = 0;
    end
  end endfunction

  function integer MAX;
    input integer LEFT, RIGHT;
  begin
    if (LEFT > RIGHT) MAX = LEFT;
    else              MAX = RIGHT;
  end endfunction

  function integer PREADDLEN;
    input integer b_len, d_len, width_d;
  begin
    if(width_d>0) PREADDLEN = MAX(b_len,d_len) + 1;
    else        PREADDLEN = b_len;
  end endfunction
  function integer PREADDMULLEN;
    input integer a_len, b_len, d_len, width_d;
  begin
    PREADDMULLEN = a_len + PREADDLEN(b_len,d_len,width_d);
  end endfunction

  localparam axb_stages = f_axb_stages(gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d);
  localparam cxd_stages = f_cxd_stages(gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d);
  localparam preadd_ab_stages = f_preadd_stages(gentype, n_inreg - axb_stages,width_b2);
  localparam preadd_cd_stages = f_preadd_stages(gentype, n_inreg - cxd_stages,width_d2);
  localparam e_stages  = (use_const>1)?n_inreg:0;
  localparam a_stages  = n_inreg - axb_stages;
  localparam b_stages  = n_inreg - axb_stages - preadd_ab_stages;
  localparam c_stages  = n_inreg - cxd_stages;
  localparam d_stages  = n_inreg - cxd_stages - preadd_cd_stages;
  localparam b2_stages  = (width_b2>0)?b_stages:0;
  localparam d2_stages  = (width_d2>0)?d_stages:0;

  localparam a_len    = width_a-signd_a+1;
  localparam b_len    = width_b-signd_b+1;
  localparam b2_len   = width_b2-signd_b2+1;
  localparam c_len    = width_c-signd_c+1;
  localparam d_len    = width_d-signd_d+1;
  localparam d2_len   = width_d2-signd_d2+1;
  localparam e_len    = width_e-signd_e+1;
  localparam bb2_len  = PREADDLEN(b_len, b2_len, width_b2);
  localparam dd2_len  = PREADDLEN(d_len, d2_len, width_d2);
  localparam axb_len  = PREADDMULLEN(a_len, b_len, b2_len, width_b2);
  localparam cxd_len  = PREADDMULLEN(c_len, d_len, d2_len, width_d2);
  localparam z_len    = width_z;

  reg [a_len-1:0]  aa  [a_stages:0];
  reg [b_len-1:0]  bb  [b_stages:0];
  reg [b2_len-1:0] bb2 [b2_stages:0];
  reg [c_len-1:0]  cc  [c_stages:0];
  reg [d_len-1:0]  dd  [d_stages:0];
  reg [d2_len-1:0] dd2 [d2_stages:0];
  reg [e_len-1:0]  ee  [e_stages:0];



  genvar i;

  // make all inputs signed
  always @(*) aa[a_stages] = signd_a ? a : {1'b0, a}; //spyglass disable W164a W164b
  always @(*) bb[b_stages] = signd_b ? b : {1'b0, b}; //spyglass disable W164a W164b
  generate if (width_b2>0) begin
    (* keep ="true" *) reg [b2_len-1:0] b2_keep;
    always @(*) b2_keep = signd_b2 ? b2 : {1'b0, b2}; //spyglass disable W164a W164b
    always @(*) bb2[b2_stages] = b2_keep;
  end endgenerate
  always @(*) cc[c_stages] = signd_c ? c : {1'b0, c}; //spyglass disable W164a W164b
  always @(*) dd[d_stages] = signd_d ? d : {1'b0, d}; //spyglass disable W164a W164b
  generate if (width_d2>0) begin
    (* keep ="true" *) reg [d2_len-1:0] d2_keep;
    always @(*) d2_keep = signd_d2 ? d2 : {1'b0, d2}; //spyglass disable W164a W164b
    always @(*) dd2[d2_stages] = d2_keep;
  end endgenerate

  generate if (use_const>0) begin
    always @(*) ee[e_stages] = signd_e ? cst : {1'b0, cst}; //spyglass disable W164a W164b

    // input registers
    if (e_stages>0) begin
    for(i = e_stages-1; i >= 0; i=i-1) begin:in_pipe_e
      if (clock_edge == 1'b1) begin:pos
        always @(posedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
      end else begin:neg
        always @(negedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
      end
    end end
  end endgenerate
  generate if (a_stages>0) begin
  for(i = a_stages-1; i >= 0; i=i-1) begin:in_pipe_a
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (b_stages>0) begin
  for(i = b_stages-1; i >= 0; i=i-1) begin:in_pipe_b
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];
    end
  end end endgenerate
  generate if (c_stages>0) begin
  for(i = c_stages-1; i >= 0; i=i-1) begin:in_pipe_c
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (d_stages>0) begin
  for(i = d_stages-1; i >= 0; i=i-1) begin:in_pipe_d
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) dd[i] <= dd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) dd[i] <= dd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (b2_stages>0) begin
  for(i = b2_stages-1; i >= 0; i=i-1) begin:in_pipe_b2
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb2[i] <= bb2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb2[i] <= bb2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (d2_stages>0) begin
  for(i = d2_stages-1; i >= 0; i=i-1) begin:in_pipe_d2
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) dd2[i] <= dd2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) dd2[i] <= dd2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg [bb2_len-1:0] b_bb2[preadd_ab_stages:0];
  reg [dd2_len-1:0] d_dd2[preadd_cd_stages:0];

  //perform first preadd
  generate
    if (width_b2>0) begin
      if (add_b2) begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]) + $signed(bb2[0]); end
      else        begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]) - $signed(bb2[0]); end
    end else      begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]); end
  endgenerate
  generate if (preadd_ab_stages>0) begin
  for(i = preadd_ab_stages-1; i >= 0; i=i-1) begin:preaddab_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) b_bb2[i] <= b_bb2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) b_bb2[i] <= b_bb2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  //perform second preadd
  generate
    if (width_d2>0) begin
      if (add_d2) begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]) + $signed(dd2[0]); end
      else        begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]) - $signed(dd2[0]); end
    end else      begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]); end
  endgenerate
  generate if (preadd_cd_stages>0) begin
  for(i = preadd_cd_stages-1; i >= 0; i=i-1) begin:preaddcd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) d_dd2[i] <= d_dd2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) d_dd2[i] <= d_dd2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // perform first multiplication
  reg [axb_len-1:0] axb[axb_stages:0];

  always @(*) axb[axb_stages] = $signed(aa[0]) * $signed(b_bb2[0]);
  generate if (axb_stages>0) begin
  for(i = axb_stages-1; i >= 0; i=i-1) begin:axb_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];
    end
  end end endgenerate

  // perform second multiplication
  reg [cxd_len-1:0] cxd[cxd_stages:0];

  always @(*) cxd[cxd_stages] = $signed(cc[0]) * $signed(d_dd2[0]);
  generate if (cxd_stages>0) begin
  for(i = cxd_stages-1; i >= 0; i=i-1) begin:cxd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cxd[i] <= cxd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cxd[i] <= cxd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg [z_len-1:0]  zz[stages-1:0];
  generate
    if (use_const>1) begin
      reg [z_len-1:0] aux_val;
      if ( isadd) begin
        always @(*) aux_val = $signed(axb[0]) + $signed(cxd[0]);
      end else begin
        always @(*) aux_val = $signed(axb[0]) - $signed(cxd[0]);
      end
      always @(*) zz[stages-1] = $signed(ee[0]) + $signed(aux_val) ;
    end else begin
      if (use_const>0) begin
        if ( isadd) begin always @(*) zz[stages-1] = $signed(axb[0]) + $signed(cxd[0]) + $signed(ee[0]); end else
                    begin always @(*) zz[stages-1] = $signed(axb[0]) - $signed(cxd[0]) + $signed(ee[0]); end
      end else begin
        if ( isadd) begin always @(*) zz[stages-1] = $signed(axb[0]) + $signed(cxd[0]); end else
                    begin always @(*) zz[stages-1] = $signed(axb[0]) - $signed(cxd[0]); end
      end
    end
  endgenerate

  // Output registers:
  generate if (stages>1) begin
  for(i = stages-2; i >= 0; i=i-1) begin:out_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // adjust output
  assign z = zz[0];
endmodule // mgc_mul2add1_pipe

//------> /cad/mentor/2024.2_1/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)
// suppress_sim_read_addr_range_errs:  0 - report errors  1 - suppress errors

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 ,
  parameter suppress_sim_read_addr_range_errs = 1 
  
)( clk,clken,d,q,radr,re,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input  re;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" , syn_ramstyle = "block" *)
  reg [data_width-1:0] mem [depth-1:0];
  integer j;
  initial for (j = 0; j < depth; j = j + 1) mem[j] = 0;
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr READ_ENABLE re
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg re_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
          re_reg <= re;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./PECore.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 03:48:28 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_PECoreRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_PECoreRun_fsm (
  clk, rst, PECoreRun_wen, fsm_output
);
  input clk;
  input rst;
  input PECoreRun_wen;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for PECore_PECore_PECoreRun_PECoreRun_fsm_1
  parameter
    PECoreRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : PECore_PECore_PECoreRun_PECoreRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // PECoreRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= PECoreRun_rlp_C_0;
    end
    else if ( PECoreRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_staller
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_staller (
  clk, rst, PECoreRun_wen, PECoreRun_wten, act_port_Push_mioi_wen_comp, rva_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PECoreRun_wen;
  output PECoreRun_wten;
  input act_port_Push_mioi_wen_comp;
  input rva_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg PECoreRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign PECoreRun_wen = act_port_Push_mioi_wen_comp & rva_out_Push_mioi_wen_comp;
  assign PECoreRun_wten = PECoreRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECoreRun_wten_reg <= 1'b0;
    end
    else begin
      PECoreRun_wten_reg <= ~ PECoreRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_wait_dp (
  weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      Datapath_for_4_ProductSum_for_acc_9_cmp_en, Datapath_for_4_ProductSum_for_acc_9_cmp_1_en,
      PECoreRun_wen, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg,
      Datapath_for_4_ProductSum_for_acc_9_cmp_cgo, Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg,
      Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_1, Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg_1
);
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output Datapath_for_4_ProductSum_for_acc_9_cmp_en;
  output Datapath_for_4_ProductSum_for_acc_9_cmp_1_en;
  input PECoreRun_wen;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg;
  input Datapath_for_4_ProductSum_for_acc_9_cmp_cgo;
  input Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg;
  input Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_1;
  input Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg_1;



  // Interconnect Declarations for Component Instantiations 
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_en = ~(PECoreRun_wen & (Datapath_for_4_ProductSum_for_acc_9_cmp_cgo
      | Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg));
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_en = ~(PECoreRun_wen & (Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_1
      | Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg_1));
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  PECoreRun_wen, rva_out_Push_mioi_oswt, rva_out_Push_mioi_biwt, rva_out_Push_mioi_bdwt,
      rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & PECoreRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt)
      & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & rva_out_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt,
      start_PopNB_mioi_biwt_pff, start_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_biwt_pff;
  input start_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & PECoreRun_wen;
  assign start_PopNB_mioi_biwt = (~ PECoreRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_biwt_pff = PECoreRun_wen & start_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp (
  clk, rst, act_port_Push_mioi_oswt, act_port_Push_mioi_wen_comp, act_port_Push_mioi_biwt,
      act_port_Push_mioi_bdwt, act_port_Push_mioi_bcwt, act_port_Push_mioi_m_data_rsc_dat,
      act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff
);
  input clk;
  input rst;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input act_port_Push_mioi_biwt;
  input act_port_Push_mioi_bdwt;
  output act_port_Push_mioi_bcwt;
  reg act_port_Push_mioi_bcwt;
  output [255:0] act_port_Push_mioi_m_data_rsc_dat;
  input [255:0] act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_wen_comp = (~ act_port_Push_mioi_oswt) | act_port_Push_mioi_biwt
      | act_port_Push_mioi_bcwt;
  assign act_port_Push_mioi_m_data_rsc_dat = {15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[240:224])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[208:192])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[176:160])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[144:128])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[112:96])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[80:64])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[48:32])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[16:0])};
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_Push_mioi_bcwt <= ~((~(act_port_Push_mioi_bcwt | act_port_Push_mioi_biwt))
          | act_port_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl (
  PECoreRun_wen, act_port_Push_mioi_oswt, act_port_Push_mioi_biwt, act_port_Push_mioi_bdwt,
      act_port_Push_mioi_bcwt, act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      act_port_Push_mioi_ccs_ccore_done_sync_vld, act_port_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_biwt;
  output act_port_Push_mioi_bdwt;
  input act_port_Push_mioi_bcwt;
  output act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input act_port_Push_mioi_ccs_ccore_done_sync_vld;
  input act_port_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_bdwt = act_port_Push_mioi_oswt & PECoreRun_wen;
  assign act_port_Push_mioi_biwt = act_port_Push_mioi_oswt & (~ act_port_Push_mioi_bcwt)
      & act_port_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & act_port_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
    (
  clk, rst, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt,
      input_port_PopNB_mioi_return_rsc_z_mxwt, input_port_PopNB_mioi_biwt, input_port_PopNB_mioi_bdwt,
      input_port_PopNB_mioi_data_data_data_rsc_z, input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_biwt;
  input input_port_PopNB_mioi_bdwt;
  input [127:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  input [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  input input_port_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg input_port_PopNB_mioi_bcwt;
  reg [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_bfwt;
  reg [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt;
  reg input_port_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_data_data_data_rsc_z_mxwt = MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z,
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt = MUX_v_8_2_2(input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z,
      input_port_PopNB_mioi_return_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      input_port_PopNB_mioi_bcwt <= ~((~(input_port_PopNB_mioi_bcwt | input_port_PopNB_mioi_biwt))
          | input_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= 8'b00000000;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( input_port_PopNB_mioi_biwt ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= input_port_PopNB_mioi_data_data_data_rsc_z;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= input_port_PopNB_mioi_data_logical_addr_rsc_z;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= input_port_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
    (
  PECoreRun_wen, PECoreRun_wten, input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_biwt,
      input_port_PopNB_mioi_bdwt, input_port_PopNB_mioi_biwt_pff, input_port_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output input_port_PopNB_mioi_biwt;
  output input_port_PopNB_mioi_bdwt;
  output input_port_PopNB_mioi_biwt_pff;
  input input_port_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_bdwt = input_port_PopNB_mioi_oswt & PECoreRun_wen;
  assign input_port_PopNB_mioi_biwt = (~ PECoreRun_wten) & input_port_PopNB_mioi_oswt;
  assign input_port_PopNB_mioi_biwt_pff = PECoreRun_wen & input_port_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [127:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  reg [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_128_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_20_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4, rva_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= 20'b00000000000000000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & PECoreRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ PECoreRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = PECoreRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, PECoreRun_wen, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_PECoreRun, rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [127:0] rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_oswt_pff(rva_out_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi (
  clk, rst, start_vld, start_rdy, start_dat, PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_vld(start_vld),
      .this_rdy(start_rdy),
      .this_dat(start_dat),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_biwt_pff(start_PopNB_mioi_biwt_iff),
      .start_PopNB_mioi_oswt_pff(start_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi (
  clk, rst, act_port_vld, act_port_rdy, act_port_dat, PECoreRun_wen, act_port_Push_mioi_oswt,
      act_port_Push_mioi_wen_comp, act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff,
      act_port_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input [255:0] act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff;
  input act_port_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_port_Push_mioi_biwt;
  wire act_port_Push_mioi_bdwt;
  wire act_port_Push_mioi_bcwt;
  wire [255:0] act_port_Push_mioi_m_data_rsc_dat;
  wire act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire act_port_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [255:0] nl_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff;
  assign nl_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff
      = {15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[240:224])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[208:192])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[176:160])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[144:128])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[112:96])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[80:64])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[48:32])
      , 15'b000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[16:0])};
  PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push  act_port_Push_mioi
      (
      .this_vld(act_port_vld),
      .this_rdy(act_port_rdy),
      .this_dat(act_port_dat),
      .m_data_rsc_dat(act_port_Push_mioi_m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt),
      .act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .act_port_Push_mioi_ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .act_port_Push_mioi_oswt_pff(act_port_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt),
      .act_port_Push_mioi_m_data_rsc_dat(act_port_Push_mioi_m_data_rsc_dat),
      .act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff(nl_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[255:0])
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi (
  clk, rst, input_port_vld, input_port_rdy, input_port_dat, PECoreRun_wen, PECoreRun_wten,
      input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt, input_port_PopNB_mioi_return_rsc_z_mxwt,
      input_port_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input input_port_vld;
  output input_port_rdy;
  input [137:0] input_port_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_port_PopNB_mioi_biwt;
  wire input_port_PopNB_mioi_bdwt;
  wire [127:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  wire input_port_PopNB_mioi_return_rsc_z;
  wire input_port_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB  input_port_PopNB_mioi
      (
      .this_vld(input_port_vld),
      .this_rdy(input_port_rdy),
      .this_dat(input_port_dat),
      .data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .return_rsc_z(input_port_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(input_port_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(input_port_PopNB_mioi_oswt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_biwt_pff(input_port_PopNB_mioi_biwt_iff),
      .input_port_PopNB_mioi_oswt_pff(input_port_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .input_port_PopNB_mioi_return_rsc_z(input_port_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt,
      rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG, weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d, Datapath_for_4_ProductSum_for_acc_9_cmp_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_c, Datapath_for_4_ProductSum_for_acc_9_cmp_en,
      Datapath_for_4_ProductSum_for_acc_9_cmp_z, Datapath_for_4_ProductSum_for_acc_9_cmp_1_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_1_c, Datapath_for_4_ProductSum_for_acc_9_cmp_1_en,
      Datapath_for_4_ProductSum_for_acc_9_cmp_1_z, Datapath_for_4_ProductSum_for_acc_9_cmp_2_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_2_c, Datapath_for_4_ProductSum_for_acc_9_cmp_2_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_3_a, Datapath_for_4_ProductSum_for_acc_9_cmp_3_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_3_z, Datapath_for_4_ProductSum_for_acc_9_cmp_4_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_4_c, Datapath_for_4_ProductSum_for_acc_9_cmp_4_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_5_a, Datapath_for_4_ProductSum_for_acc_9_cmp_5_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_5_z, Datapath_for_4_ProductSum_for_acc_9_cmp_6_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_6_c, Datapath_for_4_ProductSum_for_acc_9_cmp_6_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_7_a, Datapath_for_4_ProductSum_for_acc_9_cmp_7_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_7_z, Datapath_for_4_ProductSum_for_acc_9_cmp_8_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_8_c, Datapath_for_4_ProductSum_for_acc_9_cmp_8_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_9_a, Datapath_for_4_ProductSum_for_acc_9_cmp_9_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_9_z, Datapath_for_4_ProductSum_for_acc_9_cmp_10_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_10_c, Datapath_for_4_ProductSum_for_acc_9_cmp_10_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_11_a, Datapath_for_4_ProductSum_for_acc_9_cmp_11_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_11_z, Datapath_for_4_ProductSum_for_acc_9_cmp_12_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_12_c, Datapath_for_4_ProductSum_for_acc_9_cmp_12_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_13_a, Datapath_for_4_ProductSum_for_acc_9_cmp_13_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_13_z, Datapath_for_4_ProductSum_for_acc_9_cmp_14_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_14_c, Datapath_for_4_ProductSum_for_acc_9_cmp_14_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_15_a, Datapath_for_4_ProductSum_for_acc_9_cmp_15_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_15_z, Datapath_for_4_ProductSum_for_acc_9_cmp_16_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_16_c, Datapath_for_4_ProductSum_for_acc_9_cmp_16_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_17_a, Datapath_for_4_ProductSum_for_acc_9_cmp_17_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_17_z, Datapath_for_4_ProductSum_for_acc_9_cmp_18_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_18_c, Datapath_for_4_ProductSum_for_acc_9_cmp_18_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_19_a, Datapath_for_4_ProductSum_for_acc_9_cmp_19_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_19_z, Datapath_for_4_ProductSum_for_acc_9_cmp_20_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_20_c, Datapath_for_4_ProductSum_for_acc_9_cmp_20_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_21_a, Datapath_for_4_ProductSum_for_acc_9_cmp_21_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_21_z, Datapath_for_4_ProductSum_for_acc_9_cmp_22_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_22_c, Datapath_for_4_ProductSum_for_acc_9_cmp_22_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_23_a, Datapath_for_4_ProductSum_for_acc_9_cmp_23_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_23_z, Datapath_for_4_ProductSum_for_acc_9_cmp_24_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_24_c, Datapath_for_4_ProductSum_for_acc_9_cmp_24_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_25_a, Datapath_for_4_ProductSum_for_acc_9_cmp_25_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_25_z, Datapath_for_4_ProductSum_for_acc_9_cmp_26_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_26_c, Datapath_for_4_ProductSum_for_acc_9_cmp_26_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_27_a, Datapath_for_4_ProductSum_for_acc_9_cmp_27_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_27_z, Datapath_for_4_ProductSum_for_acc_9_cmp_28_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_28_c, Datapath_for_4_ProductSum_for_acc_9_cmp_28_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_29_a, Datapath_for_4_ProductSum_for_acc_9_cmp_29_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_29_z, Datapath_for_4_ProductSum_for_acc_9_cmp_30_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_30_c, Datapath_for_4_ProductSum_for_acc_9_cmp_30_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_31_a, Datapath_for_4_ProductSum_for_acc_9_cmp_31_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_31_z, Datapath_for_4_ProductSum_for_acc_9_cmp_32_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_32_c, Datapath_for_4_ProductSum_for_acc_9_cmp_32_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_33_a, Datapath_for_4_ProductSum_for_acc_9_cmp_33_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_33_z, Datapath_for_4_ProductSum_for_acc_9_cmp_34_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_34_c, Datapath_for_4_ProductSum_for_acc_9_cmp_34_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_35_a, Datapath_for_4_ProductSum_for_acc_9_cmp_35_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_35_z, Datapath_for_4_ProductSum_for_acc_9_cmp_36_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_36_c, Datapath_for_4_ProductSum_for_acc_9_cmp_36_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_37_a, Datapath_for_4_ProductSum_for_acc_9_cmp_37_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_37_z, Datapath_for_4_ProductSum_for_acc_9_cmp_38_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_38_c, Datapath_for_4_ProductSum_for_acc_9_cmp_38_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_39_a, Datapath_for_4_ProductSum_for_acc_9_cmp_39_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_39_z, Datapath_for_4_ProductSum_for_acc_9_cmp_40_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_40_c, Datapath_for_4_ProductSum_for_acc_9_cmp_40_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_41_a, Datapath_for_4_ProductSum_for_acc_9_cmp_41_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_41_z, Datapath_for_4_ProductSum_for_acc_9_cmp_42_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_42_c, Datapath_for_4_ProductSum_for_acc_9_cmp_42_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_43_a, Datapath_for_4_ProductSum_for_acc_9_cmp_43_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_43_z, Datapath_for_4_ProductSum_for_acc_9_cmp_44_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_44_c, Datapath_for_4_ProductSum_for_acc_9_cmp_44_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_45_a, Datapath_for_4_ProductSum_for_acc_9_cmp_45_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_45_z, Datapath_for_4_ProductSum_for_acc_9_cmp_46_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_46_c, Datapath_for_4_ProductSum_for_acc_9_cmp_46_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_47_a, Datapath_for_4_ProductSum_for_acc_9_cmp_47_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_47_z, Datapath_for_4_ProductSum_for_acc_9_cmp_48_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_48_c, Datapath_for_4_ProductSum_for_acc_9_cmp_48_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_49_a, Datapath_for_4_ProductSum_for_acc_9_cmp_49_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_49_z, Datapath_for_4_ProductSum_for_acc_9_cmp_50_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_50_c, Datapath_for_4_ProductSum_for_acc_9_cmp_50_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_51_a, Datapath_for_4_ProductSum_for_acc_9_cmp_51_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_51_z, Datapath_for_4_ProductSum_for_acc_9_cmp_52_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_52_c, Datapath_for_4_ProductSum_for_acc_9_cmp_52_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_53_a, Datapath_for_4_ProductSum_for_acc_9_cmp_53_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_53_z, Datapath_for_4_ProductSum_for_acc_9_cmp_54_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_54_c, Datapath_for_4_ProductSum_for_acc_9_cmp_54_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_55_a, Datapath_for_4_ProductSum_for_acc_9_cmp_55_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_55_z, Datapath_for_4_ProductSum_for_acc_9_cmp_56_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_56_c, Datapath_for_4_ProductSum_for_acc_9_cmp_56_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_57_a, Datapath_for_4_ProductSum_for_acc_9_cmp_57_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_57_z, Datapath_for_4_ProductSum_for_acc_9_cmp_58_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_58_c, Datapath_for_4_ProductSum_for_acc_9_cmp_58_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_59_a, Datapath_for_4_ProductSum_for_acc_9_cmp_59_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_59_z, Datapath_for_4_ProductSum_for_acc_9_cmp_60_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_60_c, Datapath_for_4_ProductSum_for_acc_9_cmp_60_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_61_a, Datapath_for_4_ProductSum_for_acc_9_cmp_61_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_61_z, Datapath_for_4_ProductSum_for_acc_9_cmp_62_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_62_c, Datapath_for_4_ProductSum_for_acc_9_cmp_62_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_63_a, Datapath_for_4_ProductSum_for_acc_9_cmp_63_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_63_z, Datapath_for_4_ProductSum_for_acc_9_cmp_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_41_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_41_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_42_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_42_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_43_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_43_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_44_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_44_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_45_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_45_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_46_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_46_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_47_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_47_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff, weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [137:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_c;
  output Datapath_for_4_ProductSum_for_acc_9_cmp_en;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_c;
  output Datapath_for_4_ProductSum_for_acc_9_cmp_1_en;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff;


  // Interconnect Declarations
  wire PECoreRun_wen;
  wire PECoreRun_wten;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  wire input_port_PopNB_mioi_return_rsc_z_mxwt;
  wire act_port_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
  wire fsm_output;
  wire pe_config_UpdateManagerCounter_if_if_unequal_tmp;
  wire [7:0] weight_mem_write_arbxbar_xbar_for_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp;
  wire while_mux_1443_tmp;
  wire while_mux_1442_tmp;
  wire while_mux_1441_tmp;
  wire while_mux_1440_tmp;
  wire while_mux_1439_tmp;
  wire while_mux_1438_tmp;
  wire while_mux_1437_tmp;
  wire while_mux_1430_tmp;
  wire while_mux_1429_tmp;
  wire while_mux_1428_tmp;
  wire while_mux_1427_tmp;
  wire while_mux_1426_tmp;
  wire while_mux_1425_tmp;
  wire while_mux_1424_tmp;
  wire while_mux_1422_tmp;
  wire while_mux_1420_tmp;
  wire while_mux_1418_tmp;
  wire while_mux_1417_tmp;
  wire while_mux_1416_tmp;
  wire while_mux_1415_tmp;
  wire while_mux_1414_tmp;
  wire while_mux_1413_tmp;
  wire while_mux_1412_tmp;
  wire while_mux_1410_tmp;
  wire while_mux_1409_tmp;
  wire while_mux_1408_tmp;
  wire while_mux_1405_tmp;
  wire weight_mem_run_3_for_weight_mem_run_3_for_and_6_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_15_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp;
  wire while_and_40_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp;
  wire weight_mem_run_3_for_weight_mem_run_3_for_and_7_tmp;
  wire weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
  wire weight_mem_run_3_for_weight_mem_run_3_for_and_1_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  wire and_dcpl_2;
  wire and_dcpl_4;
  wire and_dcpl_5;
  wire and_dcpl_24;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_33;
  wire mux_tmp;
  wire mux_tmp_4;
  wire and_dcpl_41;
  wire not_tmp_29;
  wire and_dcpl_48;
  wire or_tmp_7;
  wire or_tmp_14;
  wire or_tmp_19;
  wire or_tmp_26;
  wire or_tmp_32;
  wire and_dcpl_83;
  wire and_dcpl_90;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_96;
  wire or_dcpl_40;
  wire and_dcpl_98;
  wire and_dcpl_100;
  wire and_dcpl_102;
  wire and_dcpl_104;
  wire and_dcpl_106;
  wire or_dcpl_75;
  wire or_dcpl_80;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_167;
  wire and_dcpl_168;
  wire and_dcpl_169;
  wire and_dcpl_170;
  wire and_dcpl_172;
  wire and_dcpl_180;
  wire and_dcpl_189;
  wire and_dcpl_190;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_195;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire and_dcpl_201;
  wire and_dcpl_202;
  wire and_dcpl_203;
  wire and_dcpl_205;
  wire and_dcpl_206;
  wire and_dcpl_208;
  wire and_dcpl_209;
  wire and_dcpl_212;
  wire and_dcpl_216;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire or_dcpl_151;
  wire and_dcpl_223;
  wire and_dcpl_226;
  wire and_dcpl_227;
  wire and_dcpl_228;
  wire and_dcpl_230;
  wire or_dcpl_160;
  wire mux_tmp_31;
  wire or_tmp_47;
  wire and_dcpl_260;
  wire or_tmp_75;
  wire or_tmp_87;
  wire nor_tmp_29;
  wire mux_tmp_84;
  wire or_tmp_104;
  wire and_dcpl_277;
  wire and_dcpl_279;
  wire and_dcpl_280;
  wire and_dcpl_281;
  wire and_dcpl_295;
  wire and_dcpl_308;
  wire and_dcpl_314;
  wire and_dcpl_321;
  wire and_dcpl_346;
  wire and_dcpl_351;
  wire and_dcpl_359;
  wire and_dcpl_370;
  wire and_dcpl_373;
  wire and_dcpl_374;
  wire and_dcpl_399;
  wire and_dcpl_403;
  wire or_tmp_115;
  wire and_dcpl_433;
  wire and_dcpl_434;
  wire and_dcpl_435;
  wire or_dcpl_201;
  wire and_dcpl_458;
  wire and_dcpl_479;
  wire and_dcpl_480;
  wire mux_tmp_110;
  wire and_dcpl_488;
  wire and_dcpl_524;
  wire and_dcpl_528;
  wire and_dcpl_534;
  wire and_tmp_1;
  wire and_dcpl_537;
  wire and_tmp_2;
  wire mux_tmp_115;
  wire and_tmp_3;
  wire or_tmp_136;
  wire and_tmp_5;
  wire and_dcpl_545;
  wire and_tmp_7;
  wire mux_tmp_126;
  wire and_tmp_8;
  wire mux_tmp_130;
  wire mux_tmp_131;
  wire mux_tmp_132;
  wire and_tmp_11;
  wire and_dcpl_561;
  wire and_dcpl_562;
  wire or_dcpl_220;
  wire or_dcpl_221;
  wire or_dcpl_227;
  wire and_dcpl_578;
  wire and_dcpl_580;
  wire and_dcpl_581;
  wire and_dcpl_583;
  wire or_dcpl_231;
  wire or_dcpl_233;
  wire and_dcpl_600;
  wire or_dcpl_236;
  wire and_dcpl_643;
  wire or_dcpl_237;
  wire or_dcpl_249;
  wire or_dcpl_256;
  wire or_dcpl_257;
  wire and_dcpl_655;
  wire and_dcpl_656;
  wire and_dcpl_657;
  wire and_dcpl_659;
  wire and_dcpl_660;
  wire and_dcpl_661;
  wire and_dcpl_662;
  wire and_dcpl_663;
  wire and_dcpl_670;
  wire or_dcpl_284;
  wire or_dcpl_287;
  wire or_dcpl_291;
  wire nor_tmp_53;
  wire or_tmp_172;
  wire mux_tmp_160;
  wire nor_tmp_55;
  wire mux_tmp_161;
  wire mux_tmp_166;
  wire nand_tmp_7;
  wire mux_tmp_172;
  wire not_tmp_404;
  wire or_tmp_187;
  wire or_tmp_190;
  wire mux_tmp_180;
  wire or_tmp_193;
  wire mux_tmp_181;
  wire mux_tmp_183;
  wire mux_tmp_185;
  wire or_tmp_204;
  wire or_tmp_212;
  wire mux_tmp_195;
  wire or_tmp_219;
  wire and_dcpl_698;
  wire or_tmp_225;
  wire or_tmp_227;
  wire mux_tmp_205;
  wire mux_tmp_208;
  wire mux_tmp_211;
  wire nor_tmp_109;
  wire or_tmp_232;
  wire or_tmp_237;
  wire or_tmp_240;
  wire mux_tmp_218;
  wire or_tmp_244;
  wire or_tmp_250;
  wire or_tmp_256;
  wire and_dcpl_701;
  wire or_tmp_265;
  wire or_tmp_270;
  wire or_tmp_273;
  wire mux_tmp_241;
  wire mux_tmp_244;
  wire not_tmp_417;
  wire or_tmp_287;
  wire or_tmp_300;
  wire not_tmp_419;
  wire or_tmp_311;
  wire mux_tmp_270;
  wire mux_tmp_271;
  wire mux_tmp_274;
  wire and_dcpl_703;
  wire nor_tmp_189;
  wire mux_tmp_288;
  wire or_tmp_345;
  wire or_tmp_347;
  wire or_tmp_348;
  wire or_tmp_353;
  wire mux_tmp_307;
  wire or_tmp_358;
  wire or_tmp_362;
  wire mux_tmp_312;
  wire or_tmp_367;
  wire nor_tmp_214;
  wire or_tmp_373;
  wire nor_tmp_217;
  wire or_tmp_379;
  wire and_dcpl_706;
  wire or_tmp_389;
  wire or_tmp_395;
  wire nor_tmp_230;
  wire mux_tmp_338;
  wire or_tmp_405;
  wire or_tmp_406;
  wire or_tmp_407;
  wire or_tmp_408;
  wire or_tmp_414;
  wire or_tmp_421;
  wire and_dcpl_707;
  wire and_dcpl_712;
  wire or_tmp_442;
  wire mux_tmp_366;
  wire mux_tmp_370;
  wire mux_tmp_373;
  wire or_tmp_459;
  wire or_tmp_460;
  wire or_tmp_461;
  wire or_tmp_464;
  wire not_tmp_443;
  wire or_tmp_481;
  wire or_tmp_487;
  wire and_dcpl_717;
  wire or_tmp_496;
  wire or_tmp_509;
  wire nor_tmp_317;
  wire or_tmp_511;
  wire or_tmp_513;
  wire mux_tmp_415;
  wire not_tmp_449;
  wire nor_tmp_350;
  wire or_tmp_530;
  wire or_tmp_531;
  wire or_tmp_532;
  wire or_tmp_534;
  wire or_tmp_536;
  wire or_tmp_537;
  wire or_tmp_539;
  wire or_tmp_541;
  wire or_tmp_543;
  wire or_tmp_545;
  wire or_tmp_547;
  wire or_tmp_549;
  wire mux_tmp_435;
  wire mux_tmp_440;
  wire mux_tmp_451;
  wire mux_tmp_453;
  wire and_dcpl_720;
  wire and_dcpl_722;
  wire and_dcpl_723;
  wire and_dcpl_724;
  wire or_dcpl_295;
  wire [3:0] pe_config_manager_counter_sva_mx1;
  wire [4:0] operator_4_false_acc_sdt_sva_1;
  wire [5:0] nl_operator_4_false_acc_sdt_sva_1;
  reg [3:0] pe_config_num_manager_sva;
  wire state_0_sva_mx1;
  wire while_if_and_tmp_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiWrite_switch_lp_nor_tmp_1;
  reg pe_config_is_valid_sva;
  reg pe_config_is_zero_first_sva;
  reg pe_manager_zero_active_sva;
  reg pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  reg pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  reg PECore_UpdateFSM_switch_lp_and_7_itm_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
  reg PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  reg [8:0] operator_8_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_8_false_acc_sdt_sva_1;
  wire PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  wire PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1;
  reg PECore_RunFSM_switch_lp_nor_tmp_1;
  reg [1:0] state_2_1_sva;
  reg state_0_sva;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_3_mux_mx0w1;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_mx0w0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1;
  wire nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_5_mux_mx0w3;
  wire weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
  reg PECore_RunFSM_switch_lp_equal_tmp_1_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0;
  reg weight_mem_run_3_for_land_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg input_read_req_valid_lpi_1_dfm_1_10;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8;
  reg rva_in_reg_rw_sva_10;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_10;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  wire PECore_UpdateFSM_switch_lp_equal_tmp_6;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  wire PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
  wire PECore_UpdateFSM_switch_lp_nor_tmp_1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
  wire [7:0] pe_config_input_counter_sva_mx1;
  wire [8:0] operator_16_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_16_false_acc_sdt_sva_1;
  reg [7:0] pe_manager_num_input_sva;
  reg [7:0] pe_config_num_output_sva;
  wire PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8;
  reg weight_mem_run_3_for_land_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  wire PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  reg PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3;
  wire weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1;
  wire weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_127_sva_1;
  reg input_write_req_valid_lpi_1_dfm_1_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1;
  wire input_write_req_valid_lpi_1_dfm_5;
  wire input_mem_banks_write_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1;
  reg [14:0] pe_manager_base_input_sva;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1;
  reg rva_in_reg_rw_sva_5;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_4;
  wire PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3;
  reg rva_in_reg_rw_sva_st_1_10;
  reg input_read_req_valid_lpi_1_dfm_1_9;
  reg rva_in_reg_rw_sva_9;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
  reg rva_in_reg_rw_sva_st_1_9;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
  reg rva_in_reg_rw_sva_st_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
  reg while_stage_0_11;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  reg rva_in_reg_rw_sva_st_1_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  reg while_stage_0_5;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  reg while_stage_0_7;
  reg rva_in_reg_rw_sva_st_1_5;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1;
  reg while_stage_0_6;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_1;
  reg rva_in_reg_rw_sva_4;
  reg rva_in_reg_rw_sva_st_1_4;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3;
  reg while_stage_0_4;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  reg weight_mem_read_arbxbar_arbiters_next_7_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3;
  reg weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3;
  reg while_stage_0_3;
  reg PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  reg while_stage_0_10;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1;
  reg rva_in_reg_rw_sva_st_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_3_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_4_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_1_1_sva;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
  reg rva_in_reg_rw_sva_st_8;
  reg rva_in_reg_rw_sva_st_1_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  reg input_read_req_valid_lpi_1_dfm_1_8;
  reg rva_in_reg_rw_sva_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
  reg rva_in_reg_rw_sva_st_1_7;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  reg rva_in_reg_rw_sva_st_7;
  reg input_read_req_valid_lpi_1_dfm_1_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
  reg rva_in_reg_rw_sva_7;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
  reg rva_in_reg_rw_sva_st_6;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
  reg input_read_req_valid_lpi_1_dfm_1_6;
  reg rva_in_reg_rw_sva_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
  reg while_stage_0_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
  reg rva_in_reg_rw_sva_st_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
  reg rva_in_reg_rw_sva_st_3;
  reg rva_in_reg_rw_sva_3;
  reg input_read_req_valid_lpi_1_dfm_1_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
  reg input_read_req_valid_lpi_1_dfm_1_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
  reg input_read_req_valid_lpi_1_dfm_1_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1;
  reg [3:0] while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1;
  reg while_stage_0_9;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
  reg [1:0] state_2_1_sva_dfm_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10;
  reg while_stage_0_12;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_3;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_9;
  reg while_and_1263_itm_1;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_2;
  reg [7:0] weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs;
  wire operator_7_false_1_operator_7_false_1_or_mdf_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_3_2_0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_2_2_0;
  reg [14:0] weight_read_addrs_7_lpi_1_dfm_1;
  reg [14:0] pe_manager_base_weight_sva;
  reg [14:0] weight_read_addrs_5_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_3_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_1_lpi_1_dfm_1;
  wire [3:0] pe_manager_base_weight_sva_mx1_3_0;
  wire pe_manager_base_weight_sva_mx3_0;
  wire [14:0] pe_manager_base_weight_sva_mx2;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  wire [11:0] nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_2;
  reg [7:0] while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4;
  wire [7:0] input_write_addrs_lpi_1_dfm_2;
  wire PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
  wire Arbiter_8U_Roundrobin_pick_1_mux_429_mx1w1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_1_mux_428_mx1w1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1;
  wire while_and_221_rgt;
  wire while_and_225_rgt;
  wire while_and_229_rgt;
  wire while_and_233_rgt;
  wire while_and_237_rgt;
  wire while_and_241_rgt;
  wire while_and_245_rgt;
  wire while_and_249_rgt;
  wire while_and_253_rgt;
  wire while_and_257_rgt;
  wire while_and_261_rgt;
  wire while_and_265_rgt;
  wire while_and_269_rgt;
  wire while_and_273_rgt;
  wire while_and_277_rgt;
  wire while_and_281_rgt;
  wire while_and_285_rgt;
  wire while_and_289_rgt;
  wire while_and_293_rgt;
  wire while_and_297_rgt;
  wire while_and_301_rgt;
  wire while_and_305_rgt;
  wire while_and_309_rgt;
  wire while_and_313_rgt;
  wire while_and_317_rgt;
  wire while_and_321_rgt;
  wire while_and_325_rgt;
  wire while_and_329_rgt;
  wire while_and_333_rgt;
  wire while_and_337_rgt;
  wire while_and_341_rgt;
  wire while_and_345_rgt;
  wire while_and_349_rgt;
  wire while_and_353_rgt;
  wire while_and_357_rgt;
  wire while_and_361_rgt;
  wire while_and_365_rgt;
  wire while_and_369_rgt;
  wire while_and_373_rgt;
  wire while_and_377_rgt;
  wire while_and_381_rgt;
  wire while_and_385_rgt;
  wire while_and_389_rgt;
  wire while_and_393_rgt;
  wire while_and_397_rgt;
  wire while_and_401_rgt;
  wire while_and_405_rgt;
  wire while_and_409_rgt;
  wire while_and_413_rgt;
  wire while_and_417_rgt;
  wire while_and_421_rgt;
  wire while_and_425_rgt;
  wire while_and_429_rgt;
  wire while_and_433_rgt;
  wire while_and_437_rgt;
  wire while_and_441_rgt;
  wire while_and_445_rgt;
  wire while_and_449_rgt;
  wire while_and_453_rgt;
  wire while_and_457_rgt;
  wire while_and_461_rgt;
  wire while_and_465_rgt;
  wire while_and_469_rgt;
  wire while_and_473_rgt;
  wire while_and_477_rgt;
  wire while_and_481_rgt;
  wire while_and_485_rgt;
  wire while_and_489_rgt;
  wire while_and_493_rgt;
  wire while_and_497_rgt;
  wire while_and_501_rgt;
  wire while_and_505_rgt;
  wire while_and_509_rgt;
  wire while_and_513_rgt;
  wire while_and_517_rgt;
  wire while_and_521_rgt;
  wire while_and_525_rgt;
  wire while_and_529_rgt;
  wire while_and_533_rgt;
  wire while_and_537_rgt;
  wire while_and_541_rgt;
  wire while_and_545_rgt;
  wire while_and_549_rgt;
  wire while_and_553_rgt;
  wire while_and_557_rgt;
  wire while_and_561_rgt;
  wire while_and_565_rgt;
  wire while_and_569_rgt;
  wire while_and_573_rgt;
  wire while_and_577_rgt;
  wire while_and_581_rgt;
  wire while_and_585_rgt;
  wire while_and_589_rgt;
  wire while_and_593_rgt;
  wire while_and_597_rgt;
  wire while_and_601_rgt;
  wire while_and_605_rgt;
  wire while_and_609_rgt;
  wire while_and_613_rgt;
  wire while_and_617_rgt;
  wire while_and_621_rgt;
  wire while_and_625_rgt;
  wire while_and_629_rgt;
  wire while_and_633_rgt;
  wire while_and_637_rgt;
  wire while_and_641_rgt;
  wire while_and_645_rgt;
  wire while_and_649_rgt;
  wire while_and_653_rgt;
  wire while_and_657_rgt;
  wire while_and_661_rgt;
  wire while_and_665_rgt;
  wire while_and_669_rgt;
  wire while_and_673_rgt;
  wire while_and_677_rgt;
  wire while_and_681_rgt;
  wire while_and_685_rgt;
  wire while_and_689_rgt;
  wire while_and_693_rgt;
  wire while_and_697_rgt;
  wire while_and_701_rgt;
  wire while_and_705_rgt;
  wire while_and_709_rgt;
  wire while_and_713_rgt;
  wire while_and_717_rgt;
  wire while_and_721_rgt;
  wire while_and_725_rgt;
  wire while_and_729_rgt;
  wire while_and_733_rgt;
  wire while_and_737_rgt;
  wire while_and_741_rgt;
  wire while_and_745_rgt;
  wire while_and_749_rgt;
  wire while_and_753_rgt;
  wire while_and_757_rgt;
  wire while_and_761_rgt;
  wire while_and_765_rgt;
  wire while_and_769_rgt;
  wire while_and_773_rgt;
  wire while_and_777_rgt;
  wire while_and_781_rgt;
  wire while_and_785_rgt;
  wire while_and_789_rgt;
  wire while_and_793_rgt;
  wire while_and_797_rgt;
  wire while_and_801_rgt;
  wire while_and_805_rgt;
  wire while_and_809_rgt;
  wire while_and_813_rgt;
  wire while_and_817_rgt;
  wire while_and_821_rgt;
  wire while_and_825_rgt;
  wire while_and_829_rgt;
  wire while_and_833_rgt;
  wire while_and_837_rgt;
  wire while_and_841_rgt;
  wire while_and_845_rgt;
  wire while_and_849_rgt;
  wire while_and_853_rgt;
  wire while_and_857_rgt;
  wire while_and_861_rgt;
  wire while_and_865_rgt;
  wire while_and_869_rgt;
  wire while_and_873_rgt;
  wire while_and_877_rgt;
  wire while_and_881_rgt;
  wire while_and_885_rgt;
  wire while_and_889_rgt;
  wire while_and_893_rgt;
  wire while_and_897_rgt;
  wire while_and_901_rgt;
  wire while_and_905_rgt;
  wire while_and_909_rgt;
  wire while_and_913_rgt;
  wire while_and_917_rgt;
  wire while_and_921_rgt;
  wire while_and_925_rgt;
  wire while_and_929_rgt;
  wire while_and_933_rgt;
  wire while_and_937_rgt;
  wire while_and_941_rgt;
  wire while_and_945_rgt;
  wire while_and_949_rgt;
  wire while_and_953_rgt;
  wire while_and_957_rgt;
  wire while_and_961_rgt;
  wire while_and_965_rgt;
  wire while_and_969_rgt;
  wire while_and_973_rgt;
  wire while_and_977_rgt;
  wire while_and_981_rgt;
  wire while_and_985_rgt;
  wire while_and_989_rgt;
  wire while_and_993_rgt;
  wire while_and_997_rgt;
  wire while_and_1001_rgt;
  wire while_and_1005_rgt;
  wire while_and_1009_rgt;
  wire while_and_1013_rgt;
  wire while_and_1017_rgt;
  wire while_and_1021_rgt;
  wire while_and_1025_rgt;
  wire while_and_1029_rgt;
  wire while_and_1033_rgt;
  wire while_and_1037_rgt;
  wire while_and_1041_rgt;
  wire while_and_1045_rgt;
  wire while_and_1049_rgt;
  wire while_and_1053_rgt;
  wire while_and_1057_rgt;
  wire while_and_1061_rgt;
  wire while_and_1065_rgt;
  wire while_and_1069_rgt;
  wire while_and_1073_rgt;
  wire while_and_1077_rgt;
  wire while_and_1081_rgt;
  wire while_and_1085_rgt;
  wire while_and_1089_rgt;
  wire while_and_1093_rgt;
  wire while_and_1097_rgt;
  wire while_and_1101_rgt;
  wire while_and_1105_rgt;
  wire while_and_1109_rgt;
  wire while_and_1113_rgt;
  wire while_and_1117_rgt;
  wire while_and_1121_rgt;
  wire while_and_1125_rgt;
  wire while_and_1129_rgt;
  wire while_and_1133_rgt;
  wire while_and_1137_rgt;
  wire while_and_1141_rgt;
  wire while_and_1145_rgt;
  wire while_and_1149_rgt;
  wire while_and_1153_rgt;
  wire while_and_1157_rgt;
  wire while_and_1161_rgt;
  wire while_and_1165_rgt;
  wire while_and_1169_rgt;
  wire while_and_1173_rgt;
  wire while_and_1177_rgt;
  wire while_and_1181_rgt;
  wire while_and_1185_rgt;
  wire while_and_1189_rgt;
  wire while_and_1193_rgt;
  wire while_and_1197_rgt;
  wire while_and_1201_rgt;
  wire while_and_1205_rgt;
  wire while_and_1209_rgt;
  wire while_and_1213_rgt;
  wire while_and_1217_rgt;
  wire while_and_1221_rgt;
  wire while_and_1225_rgt;
  wire while_and_1229_rgt;
  wire while_and_1233_rgt;
  wire while_and_1237_rgt;
  wire while_and_1241_rgt;
  wire weight_mem_banks_read_1_for_mux_cse;
  wire weight_mem_banks_read_1_for_mux_1_cse;
  wire weight_mem_banks_read_1_for_mux_4_cse;
  wire weight_mem_banks_read_1_for_mux_5_cse;
  wire weight_mem_banks_read_1_for_mux_8_cse;
  wire weight_mem_banks_read_1_for_mux_9_cse;
  wire weight_mem_banks_read_1_for_mux_12_cse;
  wire weight_mem_banks_read_1_for_mux_13_cse;
  wire weight_mem_banks_read_1_for_mux_16_cse;
  wire weight_mem_banks_read_1_for_mux_17_cse;
  wire weight_mem_banks_read_1_for_mux_20_cse;
  wire weight_mem_banks_read_1_for_mux_21_cse;
  wire weight_mem_banks_read_1_for_mux_24_cse;
  wire weight_mem_banks_read_1_for_mux_25_cse;
  wire weight_mem_banks_read_1_for_mux_28_cse;
  wire weight_mem_banks_read_1_for_mux_29_cse;
  wire weight_mem_banks_write_if_for_if_mux_8_cse;
  wire weight_mem_banks_write_if_for_if_mux_9_cse;
  wire weight_mem_banks_read_for_mux_cse;
  wire weight_mem_banks_read_for_mux_1_cse;
  wire weight_mem_banks_write_if_for_if_mux_12_cse;
  wire weight_mem_banks_write_if_for_if_mux_13_cse;
  wire weight_mem_banks_read_for_mux_4_cse;
  wire weight_mem_banks_read_for_mux_5_cse;
  wire weight_mem_banks_write_if_for_if_mux_16_cse;
  wire weight_mem_banks_write_if_for_if_mux_17_cse;
  wire weight_mem_banks_read_for_mux_8_cse;
  wire weight_mem_banks_read_for_mux_9_cse;
  wire weight_mem_banks_write_if_for_if_mux_20_cse;
  wire weight_mem_banks_write_if_for_if_mux_21_cse;
  wire weight_mem_banks_read_for_mux_12_cse;
  wire weight_mem_banks_read_for_mux_13_cse;
  wire weight_mem_banks_write_if_for_if_mux_24_cse;
  wire weight_mem_banks_write_if_for_if_mux_25_cse;
  wire weight_mem_banks_read_for_mux_16_cse;
  wire weight_mem_banks_read_for_mux_17_cse;
  wire weight_mem_banks_write_if_for_if_mux_28_cse;
  wire weight_mem_banks_write_if_for_if_mux_29_cse;
  wire weight_mem_banks_read_for_mux_20_cse;
  wire weight_mem_banks_read_for_mux_21_cse;
  wire weight_mem_banks_write_if_for_if_mux_32_cse;
  wire weight_mem_banks_write_if_for_if_mux_33_cse;
  wire weight_mem_banks_read_for_mux_24_cse;
  wire weight_mem_banks_read_for_mux_25_cse;
  wire weight_mem_banks_write_if_for_if_mux_36_cse;
  wire weight_mem_banks_write_if_for_if_mux_37_cse;
  wire weight_mem_banks_read_for_mux_28_cse;
  wire weight_mem_banks_read_for_mux_29_cse;
  wire input_mem_banks_write_1_if_for_if_mux_cse;
  wire input_mem_banks_write_1_if_for_if_mux_1_cse;
  wire input_mem_banks_read_1_for_mux_cse;
  wire input_mem_banks_read_1_for_mux_1_cse;
  wire input_mem_banks_write_if_for_if_mux_cse;
  wire input_mem_banks_write_if_for_if_mux_1_cse;
  wire input_mem_banks_read_for_mux_cse;
  wire input_mem_banks_read_for_mux_1_cse;
  reg reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_63_cse;
  reg reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_56_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_act_port_Push_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire rva_out_reg_data_and_cse;
  wire weight_port_read_out_data_and_1_cse;
  wire weight_port_read_out_data_and_16_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_or_1_cse;
  wire weight_port_read_out_data_and_41_cse;
  wire weight_port_read_out_data_and_85_cse;
  reg reg_weight_mem_run_3_for_5_and_16_itm_1_cse;
  reg reg_weight_mem_run_3_for_5_and_14_itm_1_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_cse;
  reg reg_rva_in_reg_rw_sva_st_1_1_cse;
  reg [2:0] reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse;
  wire and_770_cse;
  wire and_776_cse;
  wire and_771_cse;
  wire and_766_cse;
  wire and_740_cse;
  wire and_767_cse;
  wire and_738_cse;
  wire operator_15_false_1_and_cse;
  wire pe_config_num_manager_and_cse;
  wire PECore_DecodeAxiWrite_switch_lp_and_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
  reg reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
  wire pe_manager_num_input_and_cse;
  wire or_380_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_42_cse;
  wire Arbiter_8U_Roundrobin_pick_and_37_cse;
  wire Arbiter_8U_Roundrobin_pick_or_3_cse;
  wire Arbiter_8U_Roundrobin_pick_and_7_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_30_cse;
  wire Arbiter_8U_Roundrobin_pick_and_31_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_18_cse;
  wire Arbiter_8U_Roundrobin_pick_and_25_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_8_cse;
  wire Arbiter_8U_Roundrobin_pick_and_20_cse;
  wire Arbiter_8U_Roundrobin_pick_or_1_cse;
  wire Arbiter_8U_Roundrobin_pick_and_3_cse;
  wire [1:0] state_mux_1_cse;
  wire and_319_cse;
  wire and_773_cse;
  wire and_768_cse;
  wire and_568_cse;
  wire and_803_cse;
  wire and_769_cse;
  wire and_802_cse;
  wire and_801_cse;
  wire and_666_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse;
  wire and_1114_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_3_or_cse;
  wire nand_32_cse;
  wire and_774_cse;
  wire and_804_cse;
  wire while_and_39_cse;
  wire and_162_cse;
  wire nor_404_cse;
  wire nor_405_cse;
  wire nor_412_cse;
  wire nor_409_cse;
  wire nor_410_cse;
  wire nor_413_cse;
  wire and_141_cse;
  wire and_148_cse;
  wire nor_428_cse;
  wire nor_427_cse;
  wire nor_436_cse;
  wire nand_41_cse;
  wire nand_40_cse;
  wire and_782_cse;
  wire and_797_cse;
  wire and_813_cse;
  wire and_784_cse;
  wire and_783_cse;
  wire and_817_cse;
  wire and_798_cse;
  wire and_824_cse;
  wire and_826_cse;
  wire and_825_cse;
  wire and_833_cse;
  wire and_785_cse;
  wire and_799_cse;
  wire and_800_cse;
  wire and_853_cse;
  wire and_859_cse;
  wire and_786_cse;
  wire and_787_cse;
  wire and_867_cse;
  wire and_857_cse;
  wire and_862_cse;
  wire and_858_cse;
  wire and_1100_cse;
  wire and_1101_cse;
  wire and_1092_cse;
  wire and_1094_cse;
  wire and_1093_cse;
  wire and_1095_cse;
  wire and_1098_cse;
  wire and_1097_cse;
  wire and_1096_cse;
  wire and_887_cse;
  wire and_895_cse;
  wire and_886_cse;
  wire and_1099_cse;
  wire and_906_cse;
  wire and_937_cse;
  wire and_939_cse;
  wire and_940_cse;
  wire and_938_cse;
  wire and_936_cse;
  wire and_947_cse;
  wire and_951_cse;
  wire and_789_cse;
  wire and_1107_cse;
  wire and_1110_cse;
  wire and_1108_cse;
  wire and_1106_cse;
  wire and_1109_cse;
  wire and_1111_cse;
  wire and_1118_cse;
  wire and_1009_cse;
  wire and_1008_cse;
  wire and_1119_cse;
  wire and_1024_cse;
  wire and_1034_cse;
  wire and_1028_cse;
  wire and_795_cse;
  wire and_1049_cse;
  wire and_792_cse;
  wire and_794_cse;
  wire and_793_cse;
  wire and_752_cse;
  wire and_764_cse;
  wire and_759_cse;
  wire and_758_cse;
  reg Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0;
  wire while_if_and_2_m1c;
  wire PECore_RunMac_and_cse;
  wire PECore_RunMac_and_4_cse;
  wire pe_config_is_valid_and_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_cse;
  wire Arbiter_8U_Roundrobin_pick_and_38_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_77_cse;
  wire Arbiter_8U_Roundrobin_pick_and_54_cse;
  wire and_380_cse;
  wire pe_config_input_counter_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse;
  wire and_527_cse;
  wire or_100_cse;
  wire or_79_cse;
  wire and_113_cse;
  wire and_120_cse;
  wire and_127_cse;
  wire and_134_cse;
  wire or_469_cse;
  wire or_569_cse;
  wire or_639_cse;
  wire mux_289_cse;
  wire mux_365_cse;
  wire or_811_cse;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1;
  wire PECore_DecodeAxiWrite_switch_lp_or_5_cse_1;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse;
  wire mux_285_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0;
  wire and_566_rmff;
  wire and_563_rmff;
  wire and_558_rmff;
  wire and_554_rmff;
  wire and_549_rmff;
  wire and_545_rmff;
  wire and_541_rmff;
  wire and_537_rmff;
  wire and_533_rmff;
  wire and_530_rmff;
  wire and_570_rmff;
  wire and_572_rmff;
  reg [7:0] pe_config_output_counter_sva;
  reg [7:0] pe_config_input_counter_sva;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_4_5;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4_5;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4_5;
  reg rva_out_reg_data_63_sva_dfm_4_5;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_5;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4_5;
  reg rva_out_reg_data_47_sva_dfm_4_5;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_5;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_5;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_4;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0;
  reg weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
  reg [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1;
  reg [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1;
  reg [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1;
  reg weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
  reg [7:0] weight_port_read_out_data_3_15_sva_dfm_1;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_5;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  wire [7:0] weight_port_read_out_data_0_7_sva_mx0;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  reg [7:0] weight_port_read_out_data_0_6_sva_dfm_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  reg [7:0] weight_port_read_out_data_0_9_sva_dfm_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  reg [7:0] weight_port_read_out_data_0_8_sva_dfm_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  reg [7:0] weight_port_read_out_data_0_15_sva_dfm_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
  reg [7:0] weight_port_read_out_data_6_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg [7:0] weight_port_read_out_data_6_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg [7:0] weight_port_read_out_data_6_3_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg [7:0] weight_port_read_out_data_6_2_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg [7:0] weight_port_read_out_data_6_5_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg [7:0] weight_port_read_out_data_6_4_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg [7:0] weight_port_read_out_data_6_7_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg [7:0] weight_port_read_out_data_6_6_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg [7:0] weight_port_read_out_data_6_9_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  reg [7:0] weight_port_read_out_data_6_8_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
  reg [7:0] weight_port_read_out_data_6_11_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  reg [7:0] weight_port_read_out_data_6_10_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  reg [7:0] weight_port_read_out_data_6_13_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  reg [7:0] weight_port_read_out_data_6_12_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  reg [7:0] weight_port_read_out_data_6_15_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  reg [7:0] weight_port_read_out_data_6_14_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
  reg [7:0] weight_port_read_out_data_1_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg [7:0] weight_port_read_out_data_1_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  reg [7:0] weight_port_read_out_data_1_3_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  reg [7:0] weight_port_read_out_data_1_2_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  reg [7:0] weight_port_read_out_data_1_5_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  reg [7:0] weight_port_read_out_data_1_4_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  reg [7:0] weight_port_read_out_data_1_7_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  reg [7:0] weight_port_read_out_data_1_6_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  reg [7:0] weight_port_read_out_data_1_9_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  reg [7:0] weight_port_read_out_data_1_8_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  reg [7:0] weight_port_read_out_data_1_11_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  reg [7:0] weight_port_read_out_data_1_10_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  reg [7:0] weight_port_read_out_data_1_13_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  reg [7:0] weight_port_read_out_data_1_12_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
  reg [7:0] weight_port_read_out_data_1_15_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg [7:0] weight_port_read_out_data_5_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  reg [7:0] weight_port_read_out_data_5_3_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  reg [7:0] weight_port_read_out_data_5_2_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  reg [7:0] weight_port_read_out_data_5_5_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  reg [7:0] weight_port_read_out_data_5_4_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  reg [7:0] weight_port_read_out_data_5_7_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  reg [7:0] weight_port_read_out_data_5_6_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  reg [7:0] weight_port_read_out_data_5_9_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  reg [7:0] weight_port_read_out_data_5_8_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  reg [7:0] weight_port_read_out_data_5_11_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  reg [7:0] weight_port_read_out_data_5_10_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  reg [7:0] weight_port_read_out_data_5_13_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  reg [7:0] weight_port_read_out_data_5_12_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg [7:0] weight_port_read_out_data_2_1_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  reg [7:0] weight_port_read_out_data_2_0_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  reg [7:0] weight_port_read_out_data_2_3_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  reg [7:0] weight_port_read_out_data_2_2_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  reg [7:0] weight_port_read_out_data_2_5_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  reg [7:0] weight_port_read_out_data_2_4_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  reg [7:0] weight_port_read_out_data_2_7_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  reg [7:0] weight_port_read_out_data_2_6_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  reg [7:0] weight_port_read_out_data_2_9_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  reg [7:0] weight_port_read_out_data_2_8_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  reg [7:0] weight_port_read_out_data_2_11_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  reg [7:0] weight_port_read_out_data_2_10_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  reg [7:0] weight_port_read_out_data_2_13_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  reg [7:0] weight_port_read_out_data_2_12_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
  reg [7:0] weight_port_read_out_data_2_14_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg [7:0] weight_port_read_out_data_4_1_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  reg [7:0] weight_port_read_out_data_4_0_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  reg [7:0] weight_port_read_out_data_4_3_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  reg [7:0] weight_port_read_out_data_4_2_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  reg [7:0] weight_port_read_out_data_4_5_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  reg [7:0] weight_port_read_out_data_4_4_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  reg [7:0] weight_port_read_out_data_4_7_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  reg [7:0] weight_port_read_out_data_4_6_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  reg [7:0] weight_port_read_out_data_4_9_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  reg [7:0] weight_port_read_out_data_4_8_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  reg [7:0] weight_port_read_out_data_4_11_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  reg [7:0] weight_port_read_out_data_4_10_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  reg [7:0] weight_port_read_out_data_4_13_sva_dfm_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  reg [7:0] weight_port_read_out_data_4_12_sva_dfm_1;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_4_1;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
  reg [7:0] weight_port_read_out_data_4_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
  reg [7:0] weight_port_read_out_data_3_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
  reg [7:0] weight_port_read_out_data_3_3_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
  reg [7:0] weight_port_read_out_data_3_2_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
  reg [7:0] weight_port_read_out_data_3_5_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
  reg [7:0] weight_port_read_out_data_3_4_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
  reg [7:0] weight_port_read_out_data_3_7_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
  reg [7:0] weight_port_read_out_data_3_6_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
  reg [7:0] weight_port_read_out_data_3_9_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
  reg [7:0] weight_port_read_out_data_3_8_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
  reg [7:0] weight_port_read_out_data_3_11_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
  reg [7:0] weight_port_read_out_data_3_10_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
  reg [7:0] weight_port_read_out_data_3_13_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
  reg [7:0] weight_port_read_out_data_3_12_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
  reg [7:0] weight_write_data_data_0_15_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_14_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_13_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_12_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_11_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_10_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_9_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_8_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
  reg [14:0] weight_write_addrs_lpi_1_dfm_1_2;
  reg [7:0] weight_write_data_data_0_15_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_14_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_13_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_12_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_11_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_10_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_9_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_8_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_3_2;
  reg [11:0] weight_write_addrs_lpi_1_dfm_1_3_14_3;
  reg [16:0] act_port_reg_data_240_224_sva_dfm_1_2;
  reg [16:0] act_port_reg_data_208_192_sva_dfm_1_2;
  reg [16:0] act_port_reg_data_176_160_sva_dfm_1_2;
  reg [16:0] act_port_reg_data_144_128_sva_dfm_1_1;
  reg [16:0] act_port_reg_data_112_96_sva_dfm_1_1;
  reg [16:0] act_port_reg_data_80_64_sva_dfm_1_1;
  reg [16:0] act_port_reg_data_48_32_sva_dfm_1_1;
  reg [16:0] act_port_reg_data_16_0_sva_dfm_1_2;
  wire and_dcpl;
  wire and_dcpl_725;
  wire or_dcpl;
  wire or_dcpl_296;
  wire or_dcpl_298;
  wire or_dcpl_300;
  wire or_dcpl_301;
  wire and_dcpl_737;
  wire and_676_ssc;
  wire and_677_ssc;
  wire and_678_ssc;
  wire and_680_ssc;
  wire and_683_ssc;
  wire and_686_ssc;
  reg [127:0] input_mem_banks_read_read_data_lpi_1_dfm_1_4;
  reg [127:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1;
  wire [127:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0;
  wire [119:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_5;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1;
  wire or_894_tmp;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_4;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_2;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_2;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_4;
  wire and_1147_cse;
  wire and_1148_cse;
  wire and_1149_cse;
  wire and_1150_cse;
  wire and_1151_cse;
  wire and_1152_cse;
  wire nor_626_cse;
  wire and_1156_cse;
  wire and_1157_cse;
  wire and_1158_cse;
  wire and_1159_cse;
  wire and_1160_cse;
  wire nor_627_cse;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1;
  wire [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm;
  wire mux_6_itm;
  wire mux_192_itm;
  wire mux_214_itm;
  wire mux_228_itm;
  wire mux_304_itm;
  wire mux_322_itm;
  wire mux_347_itm;
  wire mux_387_itm;
  wire mux_450_itm;
  reg weight_mem_read_arbxbar_arbiters_next_3_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_6_sva;
  reg [7:0] weight_port_read_out_data_0_7_sva;
  reg [14:0] pe_manager_base_bias_sva;
  reg pe_config_is_cluster_sva;
  reg pe_config_is_bias_sva;
  reg [3:0] pe_config_manager_counter_sva;
  reg [19:0] accum_vector_data_3_19_0_sva;
  reg [19:0] accum_vector_data_4_19_0_sva;
  reg [19:0] accum_vector_data_2_19_0_sva;
  reg [19:0] accum_vector_data_5_19_0_sva;
  reg [19:0] accum_vector_data_1_19_0_sva;
  reg [19:0] accum_vector_data_6_19_0_sva;
  reg [19:0] accum_vector_data_0_19_0_sva;
  reg [19:0] accum_vector_data_7_19_0_sva;
  reg [16:0] act_port_reg_data_112_96_sva;
  reg [16:0] act_port_reg_data_144_128_sva;
  reg [16:0] act_port_reg_data_80_64_sva;
  reg [16:0] act_port_reg_data_48_32_sva;
  reg [7:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8;
  reg [127:0] input_mem_banks_bank_a_0_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_1_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_2_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_3_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_4_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_5_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_6_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_7_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_8_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_9_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_10_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_11_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_12_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_13_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_14_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_15_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_16_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_17_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_18_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_19_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_20_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_21_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_22_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_23_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_24_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_25_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_26_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_27_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_28_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_29_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_30_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_31_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_32_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_33_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_34_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_35_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_36_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_37_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_38_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_39_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_40_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_41_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_42_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_43_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_44_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_45_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_46_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_47_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_48_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_49_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_50_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_51_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_52_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_53_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_54_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_55_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_56_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_57_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_58_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_59_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_60_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_61_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_62_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_63_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_64_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_65_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_66_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_67_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_68_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_69_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_70_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_71_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_72_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_73_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_74_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_75_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_76_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_77_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_78_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_79_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_80_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_81_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_82_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_83_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_84_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_85_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_86_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_87_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_88_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_89_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_90_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_91_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_92_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_93_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_94_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_95_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_96_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_97_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_98_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_99_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_100_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_101_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_102_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_103_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_104_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_105_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_106_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_107_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_108_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_109_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_110_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_111_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_112_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_113_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_114_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_115_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_116_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_117_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_118_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_119_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_120_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_121_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_122_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_123_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_124_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_125_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_126_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_127_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_128_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_129_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_130_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_131_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_132_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_133_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_134_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_135_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_136_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_137_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_138_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_139_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_140_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_141_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_142_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_143_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_144_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_145_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_146_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_147_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_148_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_149_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_150_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_151_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_152_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_153_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_154_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_155_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_156_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_157_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_158_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_159_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_160_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_161_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_162_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_163_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_164_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_165_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_166_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_167_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_168_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_169_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_170_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_171_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_172_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_173_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_174_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_175_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_176_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_177_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_178_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_179_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_180_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_181_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_182_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_183_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_184_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_185_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_186_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_187_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_188_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_189_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_190_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_191_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_192_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_193_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_194_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_195_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_196_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_197_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_198_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_199_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_200_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_201_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_202_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_203_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_204_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_205_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_206_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_207_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_208_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_209_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_210_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_211_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_212_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_213_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_214_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_215_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_216_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_217_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_218_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_219_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_220_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_221_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_222_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_223_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_224_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_225_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_226_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_227_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_228_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_229_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_230_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_231_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_232_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_233_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_234_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_235_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_236_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_237_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_238_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_239_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_240_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_241_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_242_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_243_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_244_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_245_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_246_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_247_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_248_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_249_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_250_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_251_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_252_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_253_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_254_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_255_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_1_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_15_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_4_15_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_15_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_1_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_8_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_9_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_10_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_11_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_12_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_13_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_14_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_15_sva_dfm_1;
  reg rva_out_reg_data_24_sva_dfm_6;
  reg rva_out_reg_data_31_sva_dfm_6;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_6;
  reg rva_out_reg_data_16_sva_dfm_6;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_6;
  reg rva_out_reg_data_8_sva_dfm_6;
  reg rva_out_reg_data_0_sva_dfm_6;
  reg [127:0] weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_6;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_6;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_6;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_6;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_6;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2;
  reg [3:0] pe_config_manager_counter_sva_dfm_3_1;
  reg [7:0] input_read_addrs_sva_1_1;
  wire [8:0] nl_input_read_addrs_sva_1_1;
  reg rva_out_reg_data_63_sva_dfm_4_4;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4_1;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4_2;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4_3;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_4_4;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4_1;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4_2;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4_3;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_4_4;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_4_2;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_4_3;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_4_4;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4_1;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4_2;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4_3;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_4_4;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_2;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_3;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_4;
  reg rva_out_reg_data_47_sva_dfm_4_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_3;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_3;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_4;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_1;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_2;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_6;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_7;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_8;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_9;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_10;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_1;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_4;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_5;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_6;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_7;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_8;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_4;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_5;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_6;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_7;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_8;
  reg [7:0] pe_config_output_counter_sva_dfm_1;
  reg [7:0] pe_config_input_counter_sva_dfm_1;
  reg [127:0] rva_in_reg_data_sva_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_8_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_9_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_10_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_11_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_12_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_13_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_14_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_15_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_2;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_1;
  reg [127:0] input_mem_banks_read_read_data_lpi_1_dfm_1_2;
  reg [127:0] input_mem_banks_read_read_data_lpi_1_dfm_1_3;
  reg [10:0] PEManager_15U_GetWeightAddr_else_acc_3_1;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
  reg [16:0] act_port_reg_data_240_224_sva_dfm_1_1;
  reg [16:0] act_port_reg_data_208_192_sva_dfm_1_1;
  reg [16:0] act_port_reg_data_176_160_sva_dfm_1_1;
  reg [16:0] act_port_reg_data_16_0_sva_dfm_1_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  reg [14:0] pe_manager_base_weight_sva_dfm_3_1;
  reg [14:0] pe_manager_base_input_sva_dfm_3_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_55_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1;
  reg [7:0] weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1;
  reg [7:0] weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_44_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1;
  reg weight_mem_run_3_for_5_and_146_itm_1;
  reg weight_mem_run_3_for_5_and_147_itm_1;
  reg weight_mem_run_3_for_5_and_148_itm_1;
  reg weight_mem_run_3_for_5_and_148_itm_2;
  reg weight_mem_run_3_for_5_and_149_itm_1;
  reg weight_mem_run_3_for_5_and_150_itm_1;
  reg weight_mem_run_3_for_5_and_150_itm_2;
  reg weight_mem_run_3_for_5_and_151_itm_1;
  reg weight_mem_run_3_for_5_and_152_itm_1;
  reg weight_mem_run_3_for_5_and_4_itm_1;
  reg weight_mem_run_3_for_5_and_6_itm_1;
  reg weight_mem_run_3_for_5_and_7_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
  reg weight_mem_run_3_for_5_and_12_itm_1;
  reg weight_mem_run_3_for_5_and_15_itm_1;
  reg weight_mem_run_3_for_5_and_100_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1;
  reg weight_mem_run_3_for_5_and_134_itm_1;
  reg weight_mem_run_3_for_5_and_134_itm_2;
  reg weight_mem_run_3_for_5_and_135_itm_1;
  reg weight_mem_run_3_for_5_and_136_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2;
  reg weight_mem_run_3_for_5_and_140_itm_1;
  reg weight_mem_run_3_for_5_and_140_itm_2;
  reg weight_mem_run_3_for_5_and_142_itm_1;
  reg weight_mem_run_3_for_5_and_143_itm_1;
  reg weight_mem_run_3_for_5_and_143_itm_2;
  reg [19:0] ProductSum_for_acc_24_itm_1;
  wire [21:0] nl_ProductSum_for_acc_24_itm_1;
  reg [18:0] ProductSum_for_acc_25_itm_1;
  wire [19:0] nl_ProductSum_for_acc_25_itm_1;
  reg [19:0] ProductSum_for_acc_40_itm_1;
  wire [21:0] nl_ProductSum_for_acc_40_itm_1;
  reg [18:0] ProductSum_for_acc_41_itm_1;
  wire [19:0] nl_ProductSum_for_acc_41_itm_1;
  reg [14:0] PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1;
  reg while_if_mux_27_itm_1;
  reg PECore_PushAxiRsp_mux_10_itm_1;
  reg PECore_PushAxiRsp_mux_23_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_9;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
  reg [119:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_8;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_3_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0;
  wire PECore_PushAxiRsp_if_else_mux_23_mx0w2;
  wire [7:0] weight_port_read_out_data_0_7_sva_dfm_mx0w2;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_33_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_20_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_19_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_18_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_17_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_15_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0;
  wire [14:0] weight_read_addrs_1_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_3_lpi_1_dfm_1_1;
  wire [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_5_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_7_lpi_1_dfm_1_1;
  wire [7:0] pe_config_output_counter_sva_mx1;
  wire pe_config_is_zero_first_sva_mx1;
  wire pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  wire [16:0] act_port_reg_data_48_32_sva_mx1;
  wire [16:0] act_port_reg_data_80_64_sva_mx1;
  wire [16:0] act_port_reg_data_112_96_sva_mx1;
  wire [16:0] act_port_reg_data_144_128_sva_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
  wire PECore_PushAxiRsp_if_else_mux_10_mx0w2;
  wire [7:0] rva_out_reg_data_127_120_sva_dfm_4_mx0w0;
  wire [7:0] rva_out_reg_data_79_72_sva_dfm_7;
  wire [7:0] rva_out_reg_data_71_64_sva_dfm_7;
  wire [7:0] rva_out_reg_data_55_48_sva_dfm_6_mx1;
  wire [6:0] rva_out_reg_data_62_56_sva_dfm_6_mx1;
  wire [6:0] rva_out_reg_data_46_40_sva_dfm_6_mx1;
  wire [3:0] rva_out_reg_data_35_32_sva_dfm_6_mx1;
  wire PECore_PushAxiRsp_mux_23_itm_1_mx0c1;
  wire [14:0] pe_manager_base_input_sva_mx2;
  wire PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  wire [7:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1;
  wire weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_4;
  wire while_and_1266_cse_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  wire PECore_UpdateFSM_switch_lp_and_2_tmp_1;
  wire [16:0] act_port_reg_data_16_0_sva_dfm_3;
  wire [16:0] act_port_reg_data_176_160_sva_dfm_3;
  wire [16:0] act_port_reg_data_208_192_sva_dfm_3;
  wire [16:0] act_port_reg_data_240_224_sva_dfm_3;
  wire rva_out_reg_data_63_sva_dfm_7;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
  wire PECore_PushAxiRsp_if_asn_79;
  wire PECore_PushAxiRsp_if_asn_81;
  wire PECore_PushAxiRsp_if_asn_83;
  wire weight_mem_run_3_for_5_asn_447;
  wire weight_mem_run_3_for_5_asn_449;
  wire weight_mem_run_3_for_5_asn_451;
  wire weight_mem_run_3_for_5_asn_453;
  wire weight_mem_run_3_for_5_asn_455;
  wire weight_mem_run_3_for_5_asn_457;
  wire weight_mem_run_3_for_5_asn_459;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420;
  wire PECore_PushAxiRsp_if_asn_87;
  wire PECore_PushAxiRsp_if_asn_89;
  wire PECore_PushAxiRsp_if_asn_91;
  wire while_asn_1039;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367;
  wire weight_mem_run_3_for_5_and_152;
  wire weight_mem_run_3_for_5_and_156;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371;
  wire [7:0] pe_manager_base_input_sva_mx1_7_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0;
  reg Datapath_for_4_ProductSum_for_acc_2_1_17;
  reg [16:0] Datapath_for_4_ProductSum_for_acc_2_1_16_0;
  reg Datapath_for_4_ProductSum_for_acc_3_1_17;
  reg [16:0] Datapath_for_4_ProductSum_for_acc_3_1_16_0;
  reg Datapath_for_2_ProductSum_for_acc_2_1_17;
  reg [16:0] Datapath_for_2_ProductSum_for_acc_2_1_16_0;
  reg Datapath_for_2_ProductSum_for_acc_3_1_17;
  reg [16:0] Datapath_for_2_ProductSum_for_acc_3_1_16_0;
  wire PECore_PushAxiRsp_if_mux1h_15;
  wire PECore_PushAxiRsp_if_mux1h_17;
  wire [7:0] weight_port_read_out_data_5_14_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_5_15_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_14_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_15_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_12_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_13_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_10_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_11_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_8_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_9_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_6_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_7_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_4_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_5_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_2_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_3_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_0_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_7_1_sva_dfm_3;
  reg reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_4_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_6_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_15_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_146_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_147_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_149_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_151_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_152_itm_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse;
  reg reg_rva_in_reg_rw_sva_2_cse;
  wire weight_mem_run_3_for_5_and_145_cse;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_7_4;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_3_0;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7_4;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_3_0;
  wire weight_mem_banks_load_store_for_else_and_68_ssc;
  reg [1:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_7_6;
  reg [5:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_5_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_6_0;
  wire weight_port_read_out_data_and_189_ssc;
  reg weight_port_read_out_data_0_0_sva_dfm_1_7;
  reg [6:0] weight_port_read_out_data_0_0_sva_dfm_1_6_0;
  wire weight_mem_banks_load_store_for_else_and_75_ssc;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1_6_0;
  wire weight_mem_banks_load_store_for_else_and_56_ssc;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1_6_0;
  wire weight_port_read_out_data_and_131_ssc;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_1_7_4;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_1_3_0;
  wire and_1155_ssc;
  reg [1:0] weight_port_read_out_data_0_2_sva_dfm_1_5_4;
  reg [3:0] weight_port_read_out_data_0_2_sva_dfm_1_3_0;
  reg weight_port_read_out_data_0_1_sva_dfm_1_7;
  reg [6:0] weight_port_read_out_data_0_1_sva_dfm_1_6_0;
  wire weight_port_read_out_data_and_185_ssc;
  reg weight_port_read_out_data_0_0_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_0_sva_dfm_2_6_0;
  wire and_1183_ssc;
  wire and_1184_ssc;
  wire and_1185_ssc;
  wire and_1186_ssc;
  wire and_1187_ssc;
  wire and_1188_ssc;
  wire nor_630_ssc;
  wire weight_port_read_out_data_0_5_sva_dfm_mx0w2_7;
  wire [6:0] weight_port_read_out_data_0_5_sva_dfm_mx0w2_6_0;
  wire and_1191_ssc;
  wire and_1193_ssc;
  wire and_1194_ssc;
  wire weight_port_read_out_data_0_4_sva_dfm_mx0w2_7;
  wire [6:0] weight_port_read_out_data_0_4_sva_dfm_mx0w2_6_0;
  wire and_1199_ssc;
  wire weight_port_read_out_data_0_0_sva_dfm_mx0w0_7;
  wire [6:0] weight_port_read_out_data_0_0_sva_dfm_mx0w0_6_0;
  reg weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
  reg [6:0] weight_port_read_out_data_0_0_sva_dfm_3_rsp_1;
  reg weight_port_read_out_data_0_1_sva_dfm_2_rsp_0;
  reg [6:0] weight_port_read_out_data_0_1_sva_dfm_2_rsp_1;
  reg [1:0] weight_port_read_out_data_0_2_sva_dfm_2_rsp_1;
  reg [3:0] weight_port_read_out_data_0_2_sva_dfm_2_rsp_2;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_2_rsp_0;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_2_rsp_1;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd;
  reg [5:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1;
  wire weight_port_read_out_data_and_182_ssc;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd;
  reg [6:0] reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1;
  reg [1:0] reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_1;
  reg [3:0] reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_2;
  reg [3:0] reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd;
  reg [3:0] reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd_1;
  wire weight_port_read_out_data_0_1_sva_mx0_7;
  wire [6:0] weight_port_read_out_data_0_1_sva_mx0_6_0;
  wire [3:0] weight_port_read_out_data_0_3_sva_mx0_7_4;
  wire [3:0] weight_port_read_out_data_0_3_sva_mx0_3_0;
  wire [1:0] weight_port_read_out_data_0_2_sva_mx0_5_4;
  wire [3:0] weight_port_read_out_data_0_2_sva_mx0_3_0;
  reg weight_port_read_out_data_0_0_sva_dfm_2_7_1;
  reg [6:0] weight_port_read_out_data_0_0_sva_dfm_2_6_0_1;
  reg weight_port_read_out_data_0_2_sva_dfm_1_1_7;
  reg weight_port_read_out_data_0_1_sva_dfm_1_1_7;
  reg [6:0] weight_port_read_out_data_0_1_sva_dfm_1_1_6_0;
  reg rva_out_reg_data_39_36_sva_dfm_4_1_3;
  reg [2:0] rva_out_reg_data_39_36_sva_dfm_4_1_2_0;
  wire weight_port_read_out_data_0_0_sva_dfm_3_7;
  wire [6:0] weight_port_read_out_data_0_0_sva_dfm_3_6_0;
  wire weight_port_read_out_data_0_5_sva_mx0_7;
  wire [6:0] weight_port_read_out_data_0_5_sva_mx0_6_0;
  wire weight_port_read_out_data_0_4_sva_mx0_7;
  wire [6:0] weight_port_read_out_data_0_4_sva_mx0_6_0;
  reg [3:0] weight_port_read_out_data_0_3_sva_7_4;
  reg [3:0] weight_port_read_out_data_0_3_sva_3_0;
  reg [1:0] weight_port_read_out_data_0_2_sva_5_4;
  reg [3:0] weight_port_read_out_data_0_2_sva_3_0;
  reg weight_port_read_out_data_0_1_sva_7;
  reg [6:0] weight_port_read_out_data_0_1_sva_6_0;
  wire weight_port_read_out_data_and_130_ssc;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_1_1_7_4;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_1_1_3_0;
  reg rva_out_reg_data_39_36_sva_dfm_4_2_3;
  reg [2:0] rva_out_reg_data_39_36_sva_dfm_4_2_2_0;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_4_7_4;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_4_3_0;
  reg [1:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_4_3;
  reg [2:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_2_0;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_6;
  reg [5:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_5_0;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_6;
  reg [5:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_5_0;
  wire rva_out_reg_data_39_36_sva_dfm_6_mx1_3;
  wire [2:0] rva_out_reg_data_39_36_sva_dfm_6_mx1_2_0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1_7;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_sva_1_7;
  wire [6:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000000;
  wire weight_port_read_out_data_0_2_sva_mx0_7;
  wire weight_port_read_out_data_0_2_sva_mx0_6;
  reg weight_port_read_out_data_0_2_sva_dfm_1_1_6;
  reg [1:0] weight_port_read_out_data_0_2_sva_dfm_1_1_5_4;
  reg [3:0] weight_port_read_out_data_0_2_sva_dfm_1_1_3_0;
  wire rva_out_reg_data_and_22_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_2_cse;
  wire rva_out_reg_data_and_25_cse;
  wire input_mem_banks_read_read_data_and_cse;
  wire weight_port_read_out_data_and_123_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_cse;
  wire act_port_reg_data_and_cse;
  wire rva_in_reg_rw_and_cse;
  wire weight_mem_run_3_for_aelse_and_cse;
  wire data_in_tmp_operator_2_for_and_1_cse;
  wire data_in_tmp_operator_2_for_and_16_cse;
  wire weight_mem_banks_read_1_read_data_and_8_cse;
  wire weight_port_read_out_data_and_136_cse;
  wire weight_mem_run_3_for_aelse_and_4_cse;
  wire weight_port_read_out_data_and_145_cse;
  wire weight_port_read_out_data_and_159_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_372_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_380_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_384_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_390_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_389_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_cse;
  wire weight_read_addrs_and_5_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_49_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_55_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_61_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_67_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_73_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_78_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_84_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_90_cse;
  wire weight_read_addrs_and_7_cse;
  wire weight_write_data_data_and_cse;
  wire weight_mem_write_arbxbar_xbar_for_1_for_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse;
  wire PECore_RunFSM_switch_lp_and_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_15_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_22_cse;
  wire Arbiter_8U_Roundrobin_pick_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_50_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_64_cse;
  wire weight_write_data_data_and_16_cse;
  wire rva_in_reg_rw_and_5_cse;
  wire PECore_UpdateFSM_switch_lp_and_9_cse;
  wire state_and_cse;
  wire PECore_PushOutput_if_and_cse;
  wire PECore_RunMac_if_and_cse;
  wire weight_mem_banks_load_store_for_else_and_1_cse;
  wire weight_mem_banks_load_store_for_else_and_cse;
  wire weight_mem_banks_load_store_for_else_and_51_cse;
  wire weight_mem_banks_load_store_for_else_and_54_cse;
  wire weight_mem_banks_load_store_for_else_and_57_cse;
  wire weight_mem_banks_load_store_for_else_and_53_cse;
  wire weight_mem_banks_load_store_for_else_and_62_cse;
  wire weight_mem_banks_load_store_for_else_and_59_cse;
  wire weight_read_addrs_and_17_cse;
  wire while_if_and_11_cse;
  wire weight_read_addrs_and_19_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse;
  wire rva_in_reg_rw_and_8_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_398_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_401_cse;
  wire weight_read_addrs_and_21_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_405_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_144_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_146_cse;
  wire weight_port_read_out_data_and_174_cse;
  wire input_mem_banks_read_read_data_and_9_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse;
  wire while_if_and_15_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_7_cse;
  wire while_if_and_6_cse;
  wire rva_out_reg_data_and_40_cse;
  wire input_read_req_valid_and_1_cse;
  wire ProductSum_for_and_cse;
  wire ProductSum_for_and_8_cse;
  wire ProductSum_for_and_2_cse;
  wire rva_in_reg_rw_and_6_cse;
  wire PECore_RunMac_if_and_1_cse;
  wire rva_in_reg_rw_and_2_cse;
  wire input_mem_banks_read_read_data_and_18_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse;
  wire pe_manager_base_weight_and_6_cse;
  wire pe_manager_base_weight_and_7_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_11_cse;
  wire while_if_and_7_cse;
  wire rva_out_reg_data_and_58_cse;
  wire input_read_req_valid_and_2_cse;
  wire PECore_RunScale_if_and_3_cse;
  wire PECore_RunMac_if_and_2_cse;
  wire rva_in_reg_rw_and_7_cse;
  wire input_mem_banks_read_read_data_and_27_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_15_cse;
  wire while_if_and_8_cse;
  wire rva_out_reg_data_and_74_cse;
  wire input_read_req_valid_and_3_cse;
  wire PECore_RunMac_if_and_3_cse;
  wire rva_in_reg_rw_and_11_cse;
  wire input_mem_banks_read_read_data_and_36_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse;
  wire PECore_RunScale_if_and_6_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_19_cse;
  wire rva_out_reg_data_and_90_cse;
  wire rva_out_reg_data_and_93_cse;
  wire rva_out_reg_data_and_98_cse;
  wire input_read_req_valid_and_4_cse;
  wire rva_out_reg_data_and_106_cse;
  wire rva_out_reg_data_and_112_cse;
  wire rva_in_reg_rw_and_3_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse;
  wire PECore_RunScale_if_and_7_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_23_cse;
  wire PECore_RunMac_if_and_6_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_24_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_27_cse;
  wire rva_out_reg_data_and_120_cse;
  wire rva_out_reg_data_and_123_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_29_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_31_cse;
  wire rva_out_reg_data_and_128_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_35_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_35_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_44_cse;
  wire while_if_and_16_cse;
  wire rva_out_reg_data_and_143_cse;
  wire rva_out_reg_data_and_111_cse;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_rsp_0;
  reg [5:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_rsp_1;
  reg [1:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_1;
  reg [2:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_2;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_5_rsp_0;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_5_rsp_1;
  reg weight_port_read_out_data_0_5_sva_rsp_0;
  reg [6:0] weight_port_read_out_data_0_5_sva_rsp_1;
  reg weight_port_read_out_data_0_4_sva_rsp_0;
  reg [6:0] weight_port_read_out_data_0_4_sva_rsp_1;
  reg rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0;
  reg [2:0] rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1;
  reg rva_out_reg_data_39_36_sva_dfm_6_rsp_0;
  reg [2:0] rva_out_reg_data_39_36_sva_dfm_6_rsp_1;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd;
  reg [2:0] reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1;
  reg reg_weight_port_read_out_data_0_2_ftd;
  reg reg_weight_port_read_out_data_0_2_ftd_1;
  reg weight_port_read_out_data_0_11_sva_dfm_2_7;
  reg weight_port_read_out_data_0_10_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_10_sva_dfm_2_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0;
  wire rva_out_reg_data_95_88_sva_dfm_7_7;
  wire rva_out_reg_data_87_80_sva_dfm_7_7;
  wire [6:0] rva_out_reg_data_87_80_sva_dfm_7_6_0;
  wire [3:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_s000000;
  wire [3:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_s000001;
  wire PECore_PushAxiRsp_if_mux1h_10_6;
  wire [5:0] PECore_PushAxiRsp_if_mux1h_10_5_0;
  wire PECore_PushAxiRsp_if_mux1h_12_6;
  wire [5:0] PECore_PushAxiRsp_if_mux1h_12_5_0;
  wire [1:0] PECore_PushAxiRsp_if_mux1h_14_4_3;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_14_2_0;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_16_5_3;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_16_2_0;
  reg weight_port_read_out_data_0_2_sva_dfm_1_7;
  reg weight_port_read_out_data_0_2_sva_dfm_1_6;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1_6;
  wire [1:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_s000000;
  wire [3:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_s000001;
  reg rva_out_reg_data_39_36_sva_dfm_4_5_3;
  reg [2:0] rva_out_reg_data_39_36_sva_dfm_4_5_2_0;
  reg [3:0] weight_port_read_out_data_0_12_sva_dfm_2_7_4;
  reg [3:0] weight_port_read_out_data_0_12_sva_dfm_2_3_0;
  reg [2:0] rva_out_reg_data_30_25_sva_dfm_6_5_3;
  reg [2:0] rva_out_reg_data_30_25_sva_dfm_6_2_0;
  reg [1:0] rva_out_reg_data_23_17_sva_dfm_6_4_3;
  reg [2:0] rva_out_reg_data_23_17_sva_dfm_6_2_0;
  reg rva_out_reg_data_15_9_sva_dfm_6_6;
  reg [5:0] rva_out_reg_data_15_9_sva_dfm_6_5_0;
  reg rva_out_reg_data_7_1_sva_dfm_6_6;
  reg [5:0] rva_out_reg_data_7_1_sva_dfm_6_5_0;
  reg rva_out_reg_data_95_88_sva_dfm_6_7;
  reg rva_out_reg_data_87_80_sva_dfm_6_7;
  reg [6:0] rva_out_reg_data_87_80_sva_dfm_6_6_0;
  reg rva_out_reg_data_87_80_sva_dfm_4_1_7;
  reg [6:0] rva_out_reg_data_87_80_sva_dfm_4_1_6_0;
  reg rva_out_reg_data_95_88_sva_dfm_4_1_7;
  wire [3:0] rva_out_reg_data_103_96_sva_dfm_4_mx0w0_7_4;
  wire [3:0] rva_out_reg_data_103_96_sva_dfm_4_mx0w0_3_0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000;
  wire [6:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000;
  wire [6:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001;
  reg weight_port_read_out_data_0_2_sva_dfm_2_rsp_0_1;
  reg weight_port_read_out_data_0_2_sva_dfm_2_rsp_0_0;
  reg weight_port_read_out_data_0_11_sva_dfm_2_6;
  reg [1:0] weight_port_read_out_data_0_11_sva_dfm_2_5_4;
  reg [3:0] weight_port_read_out_data_0_11_sva_dfm_2_3_0;
  wire rva_out_reg_data_95_88_sva_dfm_7_6;
  wire [1:0] rva_out_reg_data_95_88_sva_dfm_7_5_4;
  wire [3:0] rva_out_reg_data_95_88_sva_dfm_7_3_0;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_rsp_0;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_rsp_1;
  reg rva_out_reg_data_95_88_sva_dfm_4_2_rsp_0;
  reg rva_out_reg_data_87_80_sva_dfm_4_2_rsp_0;
  reg [6:0] rva_out_reg_data_87_80_sva_dfm_4_2_rsp_1;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_3_ftd;
  reg [6:0] reg_rva_out_reg_data_87_80_sva_dfm_4_3_ftd_1;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_1;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd;
  reg [1:0] reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd_1;
  reg [3:0] reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd_2;
  reg weight_port_read_out_data_0_13_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_13_sva_dfm_2_6_0;
  reg weight_port_read_out_data_0_14_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_14_sva_dfm_2_6_0;
  wire and_699_ssc;
  wire nor_615_ssc;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_1_7_4;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_1_3_0;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_6_7_4;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_6_3_0;
  wire rva_out_reg_data_119_112_sva_dfm_4_mx0w0_7;
  wire [6:0] rva_out_reg_data_119_112_sva_dfm_4_mx0w0_6_0;
  wire rva_out_reg_data_111_104_sva_dfm_4_mx0w0_7;
  wire [6:0] rva_out_reg_data_111_104_sva_dfm_4_mx0w0_6_0;
  wire rva_out_reg_data_87_80_sva_dfm_8_7;
  wire rva_out_reg_data_95_88_sva_dfm_8_7;
  reg rva_out_reg_data_95_88_sva_dfm_6_6;
  reg [1:0] rva_out_reg_data_95_88_sva_dfm_6_5_4;
  reg [3:0] rva_out_reg_data_95_88_sva_dfm_6_3_0;
  wire and_695_ssc;
  wire nor_613_ssc;
  reg rva_out_reg_data_119_112_sva_dfm_4_1_7;
  reg [6:0] rva_out_reg_data_119_112_sva_dfm_4_1_6_0;
  wire and_697_ssc;
  wire nor_614_ssc;
  reg rva_out_reg_data_111_104_sva_dfm_4_1_7;
  reg [6:0] rva_out_reg_data_111_104_sva_dfm_4_1_6_0;
  reg rva_out_reg_data_119_112_sva_dfm_6_7;
  reg [6:0] rva_out_reg_data_119_112_sva_dfm_6_6_0;
  reg rva_out_reg_data_111_104_sva_dfm_6_7;
  reg [6:0] rva_out_reg_data_111_104_sva_dfm_6_6_0;
  reg rva_out_reg_data_87_80_sva_dfm_4_4_7;
  reg [6:0] rva_out_reg_data_87_80_sva_dfm_4_4_6_0;
  reg rva_out_reg_data_95_88_sva_dfm_4_4_7;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_2_7_4;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_2_3_0;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_0_1;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_0_0;
  reg rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_6;
  reg [1:0] rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_5_4;
  reg [3:0] rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_3_0;
  wire rva_out_reg_data_95_88_sva_dfm_8_6;
  wire [1:0] rva_out_reg_data_95_88_sva_dfm_8_5_4;
  reg rva_out_reg_data_95_88_sva_dfm_4_5_rsp_0;
  reg rva_out_reg_data_87_80_sva_dfm_4_5_rsp_0;
  reg [6:0] rva_out_reg_data_87_80_sva_dfm_4_5_rsp_1;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_3_rsp_0;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_3_rsp_1;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_0;
  reg [1:0] reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_1;
  reg [3:0] reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_2;
  reg rva_out_reg_data_119_112_sva_dfm_4_2_rsp_0;
  reg [6:0] rva_out_reg_data_119_112_sva_dfm_4_2_rsp_1;
  reg rva_out_reg_data_111_104_sva_dfm_4_2_rsp_0;
  reg [6:0] rva_out_reg_data_111_104_sva_dfm_4_2_rsp_1;
  reg [3:0] reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd;
  reg [3:0] reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd_1;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd;
  reg [6:0] reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd_1;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd;
  reg [6:0] reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd_1;
  wire rva_out_reg_data_111_104_sva_dfm_7_7;
  wire rva_out_reg_data_119_112_sva_dfm_7_7;
  wire PECore_PushAxiRsp_if_mux1h_14_6;
  wire PECore_PushAxiRsp_if_mux1h_14_5;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_5_7_4;
  reg [3:0] rva_out_reg_data_103_96_sva_dfm_4_5_3_0;
  reg rva_out_reg_data_111_104_sva_dfm_4_4_7;
  reg [6:0] rva_out_reg_data_111_104_sva_dfm_4_4_6_0;
  reg rva_out_reg_data_119_112_sva_dfm_4_4_7;
  reg [6:0] rva_out_reg_data_119_112_sva_dfm_4_4_6_0;
  reg rva_out_reg_data_23_17_sva_dfm_6_6;
  reg rva_out_reg_data_23_17_sva_dfm_6_5;
  reg rva_out_reg_data_95_88_sva_dfm_4_4_6;
  reg [1:0] rva_out_reg_data_95_88_sva_dfm_4_4_5_4;
  reg [3:0] rva_out_reg_data_95_88_sva_dfm_4_4_3_0;
  reg rva_out_reg_data_119_112_sva_dfm_4_5_rsp_0;
  reg [6:0] rva_out_reg_data_119_112_sva_dfm_4_5_rsp_1;
  reg rva_out_reg_data_111_104_sva_dfm_4_5_rsp_0;
  reg [6:0] rva_out_reg_data_111_104_sva_dfm_4_5_rsp_1;
  reg rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_0;
  reg [1:0] rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_1;
  reg [3:0] rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_2;
  wire or_dcpl_319;
  wire or_dcpl_323;
  wire or_dcpl_324;
  wire or_dcpl_332;
  wire or_dcpl_336;
  wire or_dcpl_337;
  wire or_tmp_586;
  wire and_dcpl_886;
  wire or_tmp_622;
  wire or_tmp_623;
  wire or_tmp_638;
  wire or_tmp_639;
  wire mux_tmp_546;
  wire mux_tmp_560;
  wire mux_tmp_567;
  wire or_306_cse;
  wire and_1224_cse;
  wire xor_1_cse;
  wire and_1249_cse;
  wire mux_517_cse;
  wire and_1324_cse;
  wire and_1374_cse;
  wire and_1393_cse;
  wire nor_12_cse;
  wire and_1446_cse;
  wire and_1464_cse;
  wire and_1476_cse;
  wire and_1489_cse;
  wire and_1506_cse;
  wire and_1526_cse;
  wire nor_721_cse;
  wire and_1341_cse;
  wire nor_681_cse;
  wire nor_690_cse;
  wire and_1462_cse;
  wire and_1619_cse;
  wire nand_88_cse;
  wire or_1106_cse;
  wire or_1105_cse;
  wire and_1624_cse;
  wire and_1625_cse;
  wire or_1128_cse;
  wire and_1641_cse;
  wire and_1254_cse;
  wire and_1244_cse;
  wire and_1274_cse;
  wire or_1109_cse;
  wire and_1415_cse;
  wire and_1285_cse;
  wire and_1280_cse;
  wire and_1578_cse;
  wire mux_565_cse;
  wire and_1562_cse;
  reg reg_rva_out_reg_data_15_9_sva_dfm_9_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_7_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_7_enexo;
  reg reg_rva_out_reg_data_127_120_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_79_72_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_71_64_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo;
  reg reg_act_port_reg_data_16_0_sva_dfm_1_1_enexo;
  reg reg_act_port_reg_data_240_224_sva_dfm_1_1_enexo;
  reg reg_act_port_reg_data_208_192_sva_dfm_1_1_enexo;
  reg reg_act_port_reg_data_176_160_sva_dfm_1_1_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1;
  reg reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo;
  reg reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  reg reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_manager_base_input_enexo;
  reg reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_config_num_output_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  reg reg_rva_in_reg_data_sva_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_127_120_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_79_72_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_71_64_sva_dfm_4_3_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo;
  reg reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_2_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_2_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_127_120_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_79_72_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_71_64_sva_dfm_4_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_127_120_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_79_72_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_71_64_sva_dfm_4_1_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2;
  reg reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_1_enexo;
  reg reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_1_enexo;
  reg reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_1_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1;
  reg reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo;
  reg reg_pe_config_input_counter_sva_dfm_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo_1;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_1_2_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_1_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_1_1_enexo;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_1_enexo;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_1_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_4_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_4_1_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_3_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_3_1_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_4_1_enexo;
  reg reg_rva_out_reg_data_87_80_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_2_3_enexo;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_1_3_enexo;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_4_1_enexo;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_4_1_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_103_96_sva_dfm_4_4_1_enexo;
  reg reg_rva_out_reg_data_119_112_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_111_104_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_4_3_enexo;
  reg reg_rva_out_reg_data_95_88_sva_dfm_4_3_3_enexo;
  wire rva_out_reg_data_and_147_enex5;
  wire rva_out_reg_data_and_148_enex5;
  wire rva_out_reg_data_and_149_enex5;
  wire rva_out_reg_data_and_150_enex5;
  wire rva_out_reg_data_and_151_enex5;
  wire rva_out_reg_data_and_152_enex5;
  wire rva_out_reg_data_and_153_enex5;
  wire rva_out_reg_data_and_154_enex5;
  wire rva_out_reg_data_and_155_enex5;
  wire rva_out_reg_data_and_156_enex5;
  wire input_mem_banks_read_read_data_and_47_enex5;
  wire input_mem_banks_read_read_data_and_48_enex5;
  wire input_mem_banks_read_read_data_and_49_enex5;
  wire input_mem_banks_read_read_data_and_50_enex5;
  wire act_port_reg_data_and_19_enex5;
  wire act_port_reg_data_and_20_enex5;
  wire act_port_reg_data_and_21_enex5;
  wire act_port_reg_data_and_22_enex5;
  wire input_mem_banks_read_1_read_data_and_enex5;
  wire weight_port_read_out_data_and_enex5;
  wire weight_port_read_out_data_and_190_enex5;
  wire weight_port_read_out_data_and_191_enex5;
  wire weight_port_read_out_data_and_192_enex5;
  wire weight_port_read_out_data_and_193_enex5;
  wire weight_port_read_out_data_and_194_enex5;
  wire weight_port_read_out_data_and_195_enex5;
  wire weight_port_read_out_data_and_196_enex5;
  wire weight_port_read_out_data_and_197_enex5;
  wire weight_port_read_out_data_and_198_enex5;
  wire weight_port_read_out_data_and_199_enex5;
  wire weight_port_read_out_data_and_200_enex5;
  wire weight_port_read_out_data_and_201_enex5;
  wire weight_port_read_out_data_and_202_enex5;
  wire weight_port_read_out_data_and_203_enex5;
  wire weight_port_read_out_data_and_204_enex5;
  wire weight_port_read_out_data_and_205_enex5;
  wire weight_port_read_out_data_and_206_enex5;
  wire weight_port_read_out_data_and_207_enex5;
  wire weight_port_read_out_data_and_208_enex5;
  wire weight_port_read_out_data_and_209_enex5;
  wire weight_port_read_out_data_and_210_enex5;
  wire weight_port_read_out_data_and_211_enex5;
  wire weight_port_read_out_data_and_212_enex5;
  wire weight_port_read_out_data_and_213_enex5;
  wire weight_port_read_out_data_and_214_enex5;
  wire weight_port_read_out_data_and_215_enex5;
  wire weight_port_read_out_data_and_216_enex5;
  wire weight_port_read_out_data_and_217_enex5;
  wire weight_port_read_out_data_and_218_enex5;
  wire weight_port_read_out_data_and_219_enex5;
  wire weight_port_read_out_data_and_31_enex5;
  wire input_mem_banks_read_1_read_data_and_1_enex5;
  wire weight_read_addrs_and_28_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5;
  wire weight_write_data_data_and_48_enex5;
  wire weight_write_data_data_and_49_enex5;
  wire weight_write_data_data_and_50_enex5;
  wire weight_write_data_data_and_51_enex5;
  wire weight_write_data_data_and_52_enex5;
  wire weight_write_data_data_and_53_enex5;
  wire weight_write_data_data_and_54_enex5;
  wire weight_write_data_data_and_55_enex5;
  wire weight_write_data_data_and_56_enex5;
  wire weight_write_data_data_and_57_enex5;
  wire weight_write_data_data_and_58_enex5;
  wire weight_write_data_data_and_59_enex5;
  wire weight_write_data_data_and_60_enex5;
  wire weight_write_data_data_and_61_enex5;
  wire weight_write_data_data_and_62_enex5;
  wire weight_write_data_data_and_63_enex5;
  wire weight_write_addrs_and_enex5;
  wire weight_write_data_data_and_64_enex5;
  wire weight_write_data_data_and_65_enex5;
  wire weight_write_data_data_and_66_enex5;
  wire weight_write_data_data_and_67_enex5;
  wire weight_write_data_data_and_68_enex5;
  wire weight_write_data_data_and_69_enex5;
  wire weight_write_data_data_and_70_enex5;
  wire weight_write_data_data_and_71_enex5;
  wire weight_write_data_data_and_72_enex5;
  wire weight_write_data_data_and_73_enex5;
  wire weight_write_data_data_and_74_enex5;
  wire weight_write_data_data_and_75_enex5;
  wire weight_write_data_data_and_76_enex5;
  wire weight_write_data_data_and_77_enex5;
  wire weight_write_data_data_and_78_enex5;
  wire weight_write_data_data_and_79_enex5;
  wire weight_write_addrs_and_2_enex5;
  wire weight_read_addrs_and_29_enex5;
  wire pe_config_UpdateManagerCounter_if_if_and_enex5;
  wire weight_read_addrs_and_30_enex5;
  wire PEManager_15U_PEManagerWrite_and_enex5;
  wire weight_port_read_out_data_and_220_enex5;
  wire input_mem_banks_read_read_data_and_51_enex5;
  wire input_mem_banks_read_read_data_and_52_enex5;
  wire input_mem_banks_read_read_data_and_53_enex5;
  wire input_mem_banks_read_read_data_and_54_enex5;
  wire input_mem_banks_read_1_read_data_and_2_enex5;
  wire rva_out_reg_data_and_157_enex5;
  wire rva_out_reg_data_and_158_enex5;
  wire rva_out_reg_data_and_159_enex5;
  wire rva_out_reg_data_and_160_enex5;
  wire rva_out_reg_data_and_161_enex5;
  wire rva_out_reg_data_and_162_enex5;
  wire rva_out_reg_data_and_163_enex5;
  wire rva_out_reg_data_and_164_enex5;
  wire rva_out_reg_data_and_165_enex5;
  wire rva_out_reg_data_and_166_enex5;
  wire rva_out_reg_data_and_167_enex5;
  wire rva_out_reg_data_and_168_enex5;
  wire weight_port_read_out_data_and_221_enex5;
  wire weight_port_read_out_data_and_222_enex5;
  wire weight_mem_write_arbxbar_xbar_for_empty_and_enex5;
  wire input_mem_banks_read_read_data_and_55_enex5;
  wire input_mem_banks_read_read_data_and_56_enex5;
  wire input_mem_banks_read_read_data_and_57_enex5;
  wire input_mem_banks_read_read_data_and_58_enex5;
  wire input_mem_banks_read_1_read_data_and_3_enex5;
  wire rva_out_reg_data_and_169_enex5;
  wire rva_out_reg_data_and_170_enex5;
  wire rva_out_reg_data_and_171_enex5;
  wire weight_port_read_out_data_and_223_enex5;
  wire weight_port_read_out_data_and_224_enex5;
  wire rva_out_reg_data_and_172_enex5;
  wire rva_out_reg_data_and_173_enex5;
  wire rva_out_reg_data_and_174_enex5;
  wire rva_out_reg_data_and_175_enex5;
  wire rva_out_reg_data_and_176_enex5;
  wire rva_out_reg_data_and_177_enex5;
  wire rva_out_reg_data_and_178_enex5;
  wire rva_out_reg_data_and_179_enex5;
  wire rva_out_reg_data_and_180_enex5;
  wire rva_out_reg_data_and_181_enex5;
  wire input_mem_banks_read_read_data_and_59_enex5;
  wire input_mem_banks_read_read_data_and_60_enex5;
  wire input_mem_banks_read_read_data_and_61_enex5;
  wire input_mem_banks_read_read_data_and_62_enex5;
  wire rva_out_reg_data_and_182_enex5;
  wire rva_out_reg_data_and_183_enex5;
  wire rva_out_reg_data_and_184_enex5;
  wire rva_out_reg_data_and_185_enex5;
  wire rva_out_reg_data_and_186_enex5;
  wire rva_out_reg_data_and_187_enex5;
  wire rva_out_reg_data_and_188_enex5;
  wire rva_out_reg_data_and_189_enex5;
  wire rva_out_reg_data_and_190_enex5;
  wire rva_out_reg_data_and_191_enex5;
  wire input_mem_banks_read_read_data_and_63_enex5;
  wire input_mem_banks_read_read_data_and_64_enex5;
  wire input_mem_banks_read_read_data_and_65_enex5;
  wire rva_out_reg_data_and_192_enex5;
  wire rva_out_reg_data_and_193_enex5;
  wire rva_out_reg_data_and_194_enex5;
  wire input_mem_banks_read_read_data_and_45_enex5;
  wire rva_out_reg_data_and_195_enex5;
  wire rva_out_reg_data_and_196_enex5;
  wire rva_out_reg_data_and_197_enex5;
  wire rva_out_reg_data_and_198_enex5;
  wire rva_out_reg_data_and_199_enex5;
  wire rva_out_reg_data_and_200_enex5;
  wire rva_out_reg_data_and_201_enex5;
  wire rva_out_reg_data_and_202_enex5;
  wire input_mem_banks_read_read_data_and_46_enex5;
  wire rva_out_reg_data_and_203_enex5;
  wire rva_out_reg_data_and_204_enex5;
  wire rva_out_reg_data_and_205_enex5;
  wire rva_out_reg_data_and_206_enex5;
  wire rva_out_reg_data_and_207_enex5;
  wire rva_out_reg_data_and_208_enex5;
  wire rva_out_reg_data_and_136_enex5;
  wire rva_out_reg_data_and_209_enex5;
  wire rva_out_reg_data_and_210_enex5;
  wire rva_out_reg_data_and_211_enex5;
  wire rva_out_reg_data_and_212_enex5;
  wire rva_out_reg_data_and_213_enex5;
  wire weight_port_read_out_data_and_225_enex5;
  wire weight_port_read_out_data_and_226_enex5;
  wire weight_port_read_out_data_and_227_enex5;
  wire weight_port_read_out_data_and_228_enex5;
  wire weight_port_read_out_data_and_229_enex5;
  wire weight_port_read_out_data_and_230_enex5;
  wire weight_port_read_out_data_and_231_enex5;
  wire weight_port_read_out_data_and_232_enex5;
  wire weight_port_read_out_data_and_233_enex5;
  wire weight_port_read_out_data_and_234_enex5;
  wire weight_port_read_out_data_and_235_enex5;
  wire weight_port_read_out_data_and_236_enex5;
  wire weight_port_read_out_data_and_237_enex5;
  wire rva_out_reg_data_and_214_enex5;
  wire rva_out_reg_data_and_215_enex5;
  wire rva_out_reg_data_and_216_enex5;
  wire rva_out_reg_data_and_217_enex5;
  wire rva_out_reg_data_and_218_enex5;
  wire rva_out_reg_data_and_219_enex5;
  wire rva_out_reg_data_and_220_enex5;
  wire rva_out_reg_data_and_221_enex5;
  wire rva_out_reg_data_and_222_enex5;
  wire rva_out_reg_data_and_223_enex5;
  wire rva_out_reg_data_and_224_enex5;
  wire rva_out_reg_data_and_225_enex5;
  wire rva_out_reg_data_and_226_enex5;
  wire rva_out_reg_data_and_227_enex5;
  wire rva_out_reg_data_and_228_enex5;
  wire rva_out_reg_data_and_229_enex5;
  wire rva_out_reg_data_and_230_enex5;
  wire rva_out_reg_data_and_231_enex5;
  wire rva_out_reg_data_and_232_enex5;
  wire data_in_tmp_operator_2_for_and_tmp;
  wire data_in_tmp_operator_2_for_and_31_tmp;
  wire pe_manager_base_input_and_tmp;
  wire rva_in_reg_data_and_tmp;
  wire input_mem_banks_read_1_read_data_and_4_tmp;
  wire input_mem_banks_read_read_data_and_44_tmp;
  wire and_1441_tmp;
  wire and_1568_tmp;
  wire rva_in_reg_rw_and_4_cse;
  wire and_1209_itm;
  wire and_809_itm;
  wire mux_292_itm;
  wire mux_290_itm;
  wire mux_342_itm;
  wire mux_340_itm;
  wire PECore_PushAxiRsp_if_else_mux_24_itm;
  wire PECore_PushAxiRsp_if_else_mux_25_itm;
  wire PECore_PushAxiRsp_if_else_mux_26_itm;
  wire mux_577_itm;
  wire mux_248_cse;
  wire and_1089_cse;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27;
  wire mux_112_nl;
  wire or_334_nl;
  wire or_333_nl;
  wire mux_114_nl;
  wire or_338_nl;
  wire or_337_nl;
  wire mux_118_nl;
  wire mux_117_nl;
  wire or_343_nl;
  wire or_342_nl;
  wire mux_122_nl;
  wire mux_121_nl;
  wire or_350_nl;
  wire or_882_nl;
  wire mux_125_nl;
  wire mux_124_nl;
  wire or_356_nl;
  wire or_355_nl;
  wire mux_129_nl;
  wire mux_128_nl;
  wire or_361_nl;
  wire or_883_nl;
  wire mux_134_nl;
  wire mux_133_nl;
  wire or_367_nl;
  wire or_366_nl;
  wire mux_137_nl;
  wire mux_136_nl;
  wire or_373_nl;
  wire or_884_nl;
  wire mux_151_nl;
  wire mux_150_nl;
  wire mux_149_nl;
  wire mux_148_nl;
  wire mux_147_nl;
  wire mux_146_nl;
  wire mux_654_nl;
  wire and_1088_nl;
  wire mux_142_nl;
  wire mux_495_nl;
  wire mux_145_nl;
  wire mux_144_nl;
  wire mux_143_nl;
  wire mux_662_nl;
  wire mux_663_nl;
  wire or_378_nl;
  wire or_377_nl;
  wire or_376_nl;
  wire or_375_nl;
  wire[27:0] PECore_RunScale_if_for_2_scaled_val_mul_1_nl;
  wire[27:0] PECore_RunScale_if_for_3_scaled_val_mul_1_nl;
  wire[27:0] PECore_RunScale_if_for_4_scaled_val_mul_1_nl;
  wire[27:0] PECore_RunScale_if_for_5_scaled_val_mul_1_nl;
  wire mux_2_nl;
  wire mux_1_nl;
  wire or_6_nl;
  wire[7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl;
  wire[7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_1_nl;
  wire mux_7_nl;
  wire mux_8_nl;
  wire or_18_nl;
  wire mux_516_nl;
  wire mux_535_nl;
  wire mux_534_nl;
  wire mux_10_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_136_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_134_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_151_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_28_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl;
  wire mux_539_nl;
  wire mux_538_nl;
  wire nor_692_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_48_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl;
  wire mux_11_nl;
  wire nor_483_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_80_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_138_nl;
  wire mux_12_nl;
  wire nor_484_nl;
  wire mux_18_nl;
  wire mux_17_nl;
  wire or_39_nl;
  wire mux_16_nl;
  wire mux_15_nl;
  wire or_38_nl;
  wire mux_14_nl;
  wire or_37_nl;
  wire or_nl;
  wire mux_13_nl;
  wire or_31_nl;
  wire or_28_nl;
  wire mux_24_nl;
  wire mux_23_nl;
  wire or_54_nl;
  wire mux_22_nl;
  wire mux_21_nl;
  wire or_53_nl;
  wire mux_20_nl;
  wire or_52_nl;
  wire or_48_nl;
  wire mux_19_nl;
  wire or_43_nl;
  wire or_40_nl;
  wire mux_25_nl;
  wire mux_541_nl;
  wire mux_540_nl;
  wire nor_693_nl;
  wire nor_694_nl;
  wire[10:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl;
  wire[3:0] PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl;
  wire and_662_nl;
  wire[3:0] operator_4_false_acc_nl;
  wire[4:0] nl_operator_4_false_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_7_nl;
  wire mux_542_nl;
  wire nor_705_nl;
  wire mux_543_nl;
  wire nand_73_nl;
  wire or_1015_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_and_1_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_mux1h_15_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_nor_8_nl;
  wire[19:0] ProductSum_for_acc_38_nl;
  wire[21:0] nl_ProductSum_for_acc_38_nl;
  wire[19:0] ProductSum_for_acc_39_nl;
  wire[21:0] nl_ProductSum_for_acc_39_nl;
  wire PECore_UpdateFSM_switch_lp_not_21_nl;
  wire[19:0] ProductSum_for_acc_30_nl;
  wire[21:0] nl_ProductSum_for_acc_30_nl;
  wire[19:0] ProductSum_for_acc_31_nl;
  wire[21:0] nl_ProductSum_for_acc_31_nl;
  wire[19:0] ProductSum_for_acc_32_nl;
  wire[21:0] nl_ProductSum_for_acc_32_nl;
  wire[18:0] ProductSum_for_acc_33_nl;
  wire[19:0] nl_ProductSum_for_acc_33_nl;
  wire PECore_UpdateFSM_switch_lp_not_36_nl;
  wire[19:0] ProductSum_for_acc_26_nl;
  wire[21:0] nl_ProductSum_for_acc_26_nl;
  wire[19:0] ProductSum_for_acc_27_nl;
  wire[21:0] nl_ProductSum_for_acc_27_nl;
  wire[19:0] ProductSum_for_acc_28_nl;
  wire[21:0] nl_ProductSum_for_acc_28_nl;
  wire[18:0] ProductSum_for_acc_29_nl;
  wire[19:0] nl_ProductSum_for_acc_29_nl;
  wire PECore_UpdateFSM_switch_lp_not_34_nl;
  wire[19:0] ProductSum_for_acc_22_nl;
  wire[21:0] nl_ProductSum_for_acc_22_nl;
  wire[19:0] ProductSum_for_acc_23_nl;
  wire[21:0] nl_ProductSum_for_acc_23_nl;
  wire PECore_UpdateFSM_switch_lp_not_35_nl;
  wire mux_29_nl;
  wire mux_549_nl;
  wire mux_548_nl;
  wire mux_547_nl;
  wire mux_546_nl;
  wire nor_715_nl;
  wire mux_545_nl;
  wire nand_68_nl;
  wire mux_544_nl;
  wire nor_716_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_234_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_249_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_174_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_189_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_204_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_219_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_250_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_175_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_190_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_205_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_220_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_251_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_176_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_191_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_206_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_221_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_252_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_177_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_192_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_207_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_222_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_253_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_178_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_193_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_208_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_223_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_254_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_179_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_194_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_209_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_224_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_240_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_255_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_180_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_195_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_210_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_225_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_241_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_181_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_196_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_211_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_226_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_242_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_257_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_182_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_197_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_212_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_227_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_243_nl;
  wire[7:0] mux1h_3_nl;
  wire and_1171_nl;
  wire and_1172_nl;
  wire and_1173_nl;
  wire not_2374_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_198_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_228_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_244_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_199_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_229_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_245_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_200_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_230_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_246_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_201_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_231_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_247_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_202_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_232_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_203_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_233_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_140_nl;
  wire mux_42_nl;
  wire mux_41_nl;
  wire mux_40_nl;
  wire or_222_nl;
  wire mux_39_nl;
  wire or_221_nl;
  wire or_220_nl;
  wire mux_43_nl;
  wire or_236_nl;
  wire or_234_nl;
  wire mux_44_nl;
  wire or_241_nl;
  wire or_239_nl;
  wire mux_61_nl;
  wire mux_60_nl;
  wire mux_59_nl;
  wire mux_58_nl;
  wire mux_57_nl;
  wire mux_56_nl;
  wire mux_55_nl;
  wire mux_54_nl;
  wire or_253_nl;
  wire or_251_nl;
  wire or_249_nl;
  wire mux_53_nl;
  wire mux_52_nl;
  wire mux_655_nl;
  wire mux_51_nl;
  wire mux_474_nl;
  wire mux_657_nl;
  wire mux_50_nl;
  wire mux_47_nl;
  wire mux_468_nl;
  wire mux_659_nl;
  wire mux_49_nl;
  wire mux_48_nl;
  wire mux_464_nl;
  wire mux_46_nl;
  wire mux_505_nl;
  wire or_244_nl;
  wire mux_80_nl;
  wire mux_79_nl;
  wire mux_78_nl;
  wire mux_77_nl;
  wire mux_76_nl;
  wire mux_75_nl;
  wire mux_74_nl;
  wire mux_73_nl;
  wire or_262_nl;
  wire or_261_nl;
  wire mux_72_nl;
  wire mux_71_nl;
  wire mux_656_nl;
  wire mux_70_nl;
  wire mux_63_nl;
  wire mux_658_nl;
  wire mux_69_nl;
  wire mux_64_nl;
  wire mux_470_nl;
  wire mux_660_nl;
  wire mux_68_nl;
  wire mux_65_nl;
  wire mux_466_nl;
  wire mux_472_nl;
  wire mux_661_nl;
  wire mux_67_nl;
  wire mux_66_nl;
  wire mux_476_nl;
  wire mux_477_nl;
  wire mux_478_nl;
  wire mux_506_nl;
  wire or_256_nl;
  wire mux_89_nl;
  wire or_270_nl;
  wire mux_88_nl;
  wire mux_87_nl;
  wire mux_86_nl;
  wire nor_503_nl;
  wire mux_85_nl;
  wire and_267_nl;
  wire or_266_nl;
  wire mux_93_nl;
  wire mux_92_nl;
  wire mux_91_nl;
  wire or_279_nl;
  wire or_876_nl;
  wire nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_nl;
  wire mux_90_nl;
  wire or_277_nl;
  wire nand_2_nl;
  wire nor_35_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_1_nl;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_37_nl;
  wire or_274_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl;
  wire[7:0] PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_1_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_27_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_135_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_142_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_132_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl;
  wire mux_95_nl;
  wire[27:0] PECore_RunScale_if_for_1_scaled_val_mul_1_nl;
  wire[27:0] PECore_RunScale_if_for_6_scaled_val_mul_1_nl;
  wire[27:0] PECore_RunScale_if_for_7_scaled_val_mul_1_nl;
  wire[27:0] PECore_RunScale_if_for_8_scaled_val_mul_1_nl;
  wire[16:0] act_port_reg_operator_for_act_port_reg_operator_for_and_nl;
  wire[16:0] act_port_reg_operator_for_act_port_reg_operator_for_and_1_nl;
  wire[16:0] act_port_reg_operator_for_act_port_reg_operator_for_and_2_nl;
  wire[16:0] act_port_reg_operator_for_act_port_reg_operator_for_and_3_nl;
  wire[19:0] ProductSum_for_acc_nl;
  wire[21:0] nl_ProductSum_for_acc_nl;
  wire[19:0] ProductSum_for_acc_50_nl;
  wire[21:0] nl_ProductSum_for_acc_50_nl;
  wire[19:0] ProductSum_for_acc_51_nl;
  wire[21:0] nl_ProductSum_for_acc_51_nl;
  wire[18:0] ProductSum_for_acc_52_nl;
  wire[19:0] nl_ProductSum_for_acc_52_nl;
  wire PECore_UpdateFSM_switch_lp_not_37_nl;
  wire[19:0] ProductSum_for_acc_46_nl;
  wire[21:0] nl_ProductSum_for_acc_46_nl;
  wire[19:0] ProductSum_for_acc_47_nl;
  wire[21:0] nl_ProductSum_for_acc_47_nl;
  wire[19:0] ProductSum_for_acc_48_nl;
  wire[21:0] nl_ProductSum_for_acc_48_nl;
  wire[18:0] ProductSum_for_acc_49_nl;
  wire[19:0] nl_ProductSum_for_acc_49_nl;
  wire PECore_UpdateFSM_switch_lp_not_23_nl;
  wire[19:0] ProductSum_for_acc_42_nl;
  wire[21:0] nl_ProductSum_for_acc_42_nl;
  wire[19:0] ProductSum_for_acc_43_nl;
  wire[21:0] nl_ProductSum_for_acc_43_nl;
  wire[19:0] ProductSum_for_acc_44_nl;
  wire[21:0] nl_ProductSum_for_acc_44_nl;
  wire[18:0] ProductSum_for_acc_45_nl;
  wire[19:0] nl_ProductSum_for_acc_45_nl;
  wire PECore_UpdateFSM_switch_lp_not_38_nl;
  wire[19:0] ProductSum_for_acc_34_nl;
  wire[21:0] nl_ProductSum_for_acc_34_nl;
  wire[19:0] ProductSum_for_acc_35_nl;
  wire[21:0] nl_ProductSum_for_acc_35_nl;
  wire[19:0] ProductSum_for_acc_36_nl;
  wire[21:0] nl_ProductSum_for_acc_36_nl;
  wire[18:0] ProductSum_for_acc_37_nl;
  wire[19:0] nl_ProductSum_for_acc_37_nl;
  wire PECore_UpdateFSM_switch_lp_not_39_nl;
  wire[7:0] input_mem_banks_read_1_for_mux_nl;
  wire and_1206_nl;
  wire mux_96_nl;
  wire nor_462_nl;
  wire and_693_nl;
  wire nor_612_nl;
  wire weight_port_read_out_data_mux_144_nl;
  wire and_703_nl;
  wire nor_616_nl;
  wire mux_33_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_248_nl;
  wire mux_104_nl;
  wire mux_103_nl;
  wire mux_102_nl;
  wire mux_101_nl;
  wire mux_100_nl;
  wire mux_99_nl;
  wire mux_98_nl;
  wire mux_97_nl;
  wire mux_554_nl;
  wire mux_553_nl;
  wire mux_552_nl;
  wire mux_551_nl;
  wire or_1108_nl;
  wire or_1107_nl;
  wire[14:0] while_if_while_if_and_2_nl;
  wire or_465_nl;
  wire mux_105_nl;
  wire or_317_nl;
  wire mux_107_nl;
  wire mux_106_nl;
  wire mux_108_nl;
  wire and_805_nl;
  wire mux_109_nl;
  wire nor_465_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_6_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl;
  wire[7:0] mux1h_4_nl;
  wire not_2376_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_56_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_57_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_58_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_59_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_60_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_61_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_73_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_83_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_98_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_99_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_103_nl;
  wire[14:0] PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_nl;
  wire[14:0] nl_operator_15_false_acc_nl;
  wire[14:0] PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[12:0] operator_15_false_acc_1_nl;
  wire[13:0] nl_operator_15_false_acc_1_nl;
  wire[14:0] PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_2_nl;
  wire[14:0] nl_operator_15_false_acc_2_nl;
  wire[14:0] PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl;
  wire[7:0] pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl;
  wire[7:0] operator_8_false_acc_nl;
  wire[8:0] nl_operator_8_false_acc_nl;
  wire pe_config_UpdateInputCounter_not_nl;
  wire pe_config_input_counter_nand_nl;
  wire[7:0] pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl;
  wire[7:0] operator_8_false_1_acc_nl;
  wire[8:0] nl_operator_8_false_1_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_9_nl;
  wire pe_config_output_counter_nand_nl;
  wire while_and_152_nl;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl;
  wire while_if_or_nl;
  wire while_if_and_4_nl;
  wire[16:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_nl;
  wire PECore_UpdateFSM_switch_lp_not_27_nl;
  wire[16:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_nl;
  wire PECore_UpdateFSM_switch_lp_not_28_nl;
  wire[16:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_nl;
  wire PECore_UpdateFSM_switch_lp_not_29_nl;
  wire[16:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_11_nl;
  wire PECore_UpdateFSM_switch_lp_not_19_nl;
  wire PECore_PushAxiRsp_mux_24_nl;
  wire[7:0] while_if_while_if_and_24_nl;
  wire[7:0] while_if_while_if_and_30_nl;
  wire[7:0] while_if_while_if_and_31_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_nl;
  wire weight_mem_banks_load_store_1_for_else_else_or_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_4_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_6_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_8_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_21_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_265_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_69_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_202_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_238_nl;
  wire mux_237_nl;
  wire mux_236_nl;
  wire or_566_nl;
  wire or_561_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl;
  wire while_mux_1435_nl;
  wire while_mux_1436_nl;
  wire mux_284_nl;
  wire or_628_nl;
  wire mux_283_nl;
  wire or_622_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl;
  wire mux_286_nl;
  wire nor_617_nl;
  wire nor_618_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_337_nl;
  wire mux_336_nl;
  wire mux_335_nl;
  wire mux_334_nl;
  wire or_695_nl;
  wire or_694_nl;
  wire mux_333_nl;
  wire mux_332_nl;
  wire or_693_nl;
  wire or_692_nl;
  wire mux_331_nl;
  wire or_691_nl;
  wire or_685_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl;
  wire while_mux_1421_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_608_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl;
  wire nor_621_nl;
  wire mux_362_nl;
  wire or_885_nl;
  wire or_886_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_32_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl;
  wire mux_407_nl;
  wire nor_622_nl;
  wire nor_623_nl;
  wire mux_406_nl;
  wire mux_405_nl;
  wire mux_404_nl;
  wire or_794_nl;
  wire or_793_nl;
  wire or_792_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl;
  wire PECore_UpdateFSM_switch_lp_mux1h_14_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl;
  wire PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl;
  wire PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_111_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_144_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_127_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_159_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_102_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_150_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_118_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_165_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_105_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_151_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_121_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_166_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_104_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_152_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_120_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_167_nl;
  wire PECore_UpdateFSM_switch_lp_not_31_nl;
  wire PECore_UpdateFSM_switch_lp_not_32_nl;
  wire PECore_UpdateFSM_switch_lp_not_33_nl;
  wire PECore_UpdateFSM_switch_lp_not_30_nl;
  wire[7:0] PEManager_15U_GetInputAddr_acc_nl;
  wire[8:0] nl_PEManager_15U_GetInputAddr_acc_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_589_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_590_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_591_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_592_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_593_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_594_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_601_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_602_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_603_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_604_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_605_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_606_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_607_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_609_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_611_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_612_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_613_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_614_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_615_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_616_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_618_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_619_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_622_nl;
  wire or_5_nl;
  wire or_4_nl;
  wire or_11_nl;
  wire nand_nl;
  wire mux_3_nl;
  wire or_13_nl;
  wire mux_28_nl;
  wire nor_433_nl;
  wire or_193_nl;
  wire mux_30_nl;
  wire or_209_nl;
  wire mux_83_nl;
  wire mux_82_nl;
  wire mux_81_nl;
  wire or_268_nl;
  wire mux_111_nl;
  wire or_332_nl;
  wire mux_113_nl;
  wire or_336_nl;
  wire or_341_nl;
  wire mux_116_nl;
  wire or_340_nl;
  wire mux_119_nl;
  wire and_547_nl;
  wire or_347_nl;
  wire mux_120_nl;
  wire or_346_nl;
  wire mux_123_nl;
  wire or_352_nl;
  wire or_360_nl;
  wire mux_127_nl;
  wire or_359_nl;
  wire or_363_nl;
  wire and_562_nl;
  wire and_561_nl;
  wire mux_135_nl;
  wire or_370_nl;
  wire or_466_nl;
  wire mux_165_nl;
  wire mux_164_nl;
  wire mux_163_nl;
  wire or_471_nl;
  wire mux_162_nl;
  wire or_470_nl;
  wire or_468_nl;
  wire mux_171_nl;
  wire mux_170_nl;
  wire mux_169_nl;
  wire mux_168_nl;
  wire mux_167_nl;
  wire or_475_nl;
  wire nor_551_nl;
  wire mux_178_nl;
  wire nor_552_nl;
  wire mux_177_nl;
  wire mux_176_nl;
  wire mux_175_nl;
  wire mux_174_nl;
  wire nand_8_nl;
  wire nor_553_nl;
  wire mux_173_nl;
  wire or_473_nl;
  wire or_480_nl;
  wire or_491_nl;
  wire or_493_nl;
  wire mux_182_nl;
  wire or_492_nl;
  wire or_486_nl;
  wire mux_184_nl;
  wire mux_186_nl;
  wire or_497_nl;
  wire or_494_nl;
  wire mux_191_nl;
  wire mux_190_nl;
  wire mux_189_nl;
  wire mux_188_nl;
  wire or_506_nl;
  wire mux_187_nl;
  wire or_504_nl;
  wire or_501_nl;
  wire or_500_nl;
  wire mux_194_nl;
  wire mux_193_nl;
  wire or_512_nl;
  wire or_511_nl;
  wire or_510_nl;
  wire or_509_nl;
  wire mux_201_nl;
  wire mux_200_nl;
  wire mux_199_nl;
  wire mux_198_nl;
  wire mux_197_nl;
  wire mux_196_nl;
  wire or_519_nl;
  wire or_518_nl;
  wire or_517_nl;
  wire or_516_nl;
  wire or_513_nl;
  wire mux_204_nl;
  wire mux_203_nl;
  wire or_523_nl;
  wire or_521_nl;
  wire mux_207_nl;
  wire mux_206_nl;
  wire nand_9_nl;
  wire mux_210_nl;
  wire mux_209_nl;
  wire nand_10_nl;
  wire mux_213_nl;
  wire mux_212_nl;
  wire or_525_nl;
  wire or_524_nl;
  wire mux_217_nl;
  wire mux_216_nl;
  wire mux_215_nl;
  wire or_530_nl;
  wire or_529_nl;
  wire or_528_nl;
  wire mux_221_nl;
  wire mux_220_nl;
  wire mux_219_nl;
  wire or_537_nl;
  wire or_536_nl;
  wire mux_227_nl;
  wire mux_226_nl;
  wire mux_225_nl;
  wire or_544_nl;
  wire or_543_nl;
  wire mux_224_nl;
  wire mux_223_nl;
  wire or_542_nl;
  wire or_541_nl;
  wire mux_222_nl;
  wire or_540_nl;
  wire or_533_nl;
  wire mux_235_nl;
  wire mux_234_nl;
  wire mux_233_nl;
  wire mux_232_nl;
  wire nor_555_nl;
  wire nor_556_nl;
  wire nor_557_nl;
  wire nor_558_nl;
  wire mux_231_nl;
  wire mux_230_nl;
  wire mux_229_nl;
  wire nor_559_nl;
  wire nor_560_nl;
  wire nor_561_nl;
  wire nor_562_nl;
  wire mux_240_nl;
  wire mux_239_nl;
  wire or_567_nl;
  wire mux_243_nl;
  wire mux_242_nl;
  wire or_571_nl;
  wire or_570_nl;
  wire nand_11_nl;
  wire nor_565_nl;
  wire mux_256_nl;
  wire mux_255_nl;
  wire nor_566_nl;
  wire mux_254_nl;
  wire mux_253_nl;
  wire mux_252_nl;
  wire mux_251_nl;
  wire mux_250_nl;
  wire nand_12_nl;
  wire mux_249_nl;
  wire or_576_nl;
  wire mux_262_nl;
  wire or_593_nl;
  wire or_592_nl;
  wire mux_268_nl;
  wire nor_567_nl;
  wire mux_267_nl;
  wire nor_568_nl;
  wire mux_266_nl;
  wire mux_265_nl;
  wire mux_264_nl;
  wire or_600_nl;
  wire mux_263_nl;
  wire or_598_nl;
  wire or_597_nl;
  wire or_596_nl;
  wire mux_261_nl;
  wire nor_569_nl;
  wire nor_570_nl;
  wire or_611_nl;
  wire or_610_nl;
  wire or_613_nl;
  wire mux_282_nl;
  wire mux_281_nl;
  wire mux_280_nl;
  wire or_621_nl;
  wire or_620_nl;
  wire mux_279_nl;
  wire mux_278_nl;
  wire mux_277_nl;
  wire mux_276_nl;
  wire mux_275_nl;
  wire or_618_nl;
  wire or_617_nl;
  wire or_616_nl;
  wire or_615_nl;
  wire mux_273_nl;
  wire mux_272_nl;
  wire or_612_nl;
  wire or_609_nl;
  wire or_608_nl;
  wire or_637_nl;
  wire mux_287_nl;
  wire or_636_nl;
  wire or_635_nl;
  wire nand_14_nl;
  wire nand_13_nl;
  wire mux_303_nl;
  wire mux_302_nl;
  wire mux_301_nl;
  wire mux_300_nl;
  wire mux_299_nl;
  wire mux_298_nl;
  wire mux_297_nl;
  wire mux_296_nl;
  wire mux_295_nl;
  wire mux_294_nl;
  wire mux_293_nl;
  wire mux_291_nl;
  wire mux_305_nl;
  wire mux_306_nl;
  wire or_651_nl;
  wire or_650_nl;
  wire mux_310_nl;
  wire mux_309_nl;
  wire mux_308_nl;
  wire or_652_nl;
  wire or_649_nl;
  wire mux_311_nl;
  wire or_660_nl;
  wire or_659_nl;
  wire mux_315_nl;
  wire mux_314_nl;
  wire mux_313_nl;
  wire or_661_nl;
  wire or_658_nl;
  wire mux_321_nl;
  wire mux_320_nl;
  wire mux_319_nl;
  wire or_667_nl;
  wire or_666_nl;
  wire mux_318_nl;
  wire mux_317_nl;
  wire or_665_nl;
  wire or_664_nl;
  wire mux_316_nl;
  wire or_663_nl;
  wire or_654_nl;
  wire mux_329_nl;
  wire mux_328_nl;
  wire mux_327_nl;
  wire mux_326_nl;
  wire nor_571_nl;
  wire nor_572_nl;
  wire nor_573_nl;
  wire nor_574_nl;
  wire mux_325_nl;
  wire mux_324_nl;
  wire mux_323_nl;
  wire nor_575_nl;
  wire nor_576_nl;
  wire nor_577_nl;
  wire nor_578_nl;
  wire or_699_nl;
  wire or_697_nl;
  wire nand_18_nl;
  wire nand_16_nl;
  wire mux_346_nl;
  wire mux_345_nl;
  wire mux_344_nl;
  wire mux_343_nl;
  wire mux_341_nl;
  wire mux_339_nl;
  wire mux_350_nl;
  wire mux_349_nl;
  wire mux_348_nl;
  wire or_708_nl;
  wire or_707_nl;
  wire or_706_nl;
  wire mux_353_nl;
  wire mux_352_nl;
  wire mux_351_nl;
  wire or_715_nl;
  wire or_714_nl;
  wire or_713_nl;
  wire mux_360_nl;
  wire mux_359_nl;
  wire mux_358_nl;
  wire mux_357_nl;
  wire or_721_nl;
  wire or_720_nl;
  wire mux_356_nl;
  wire mux_355_nl;
  wire or_719_nl;
  wire or_718_nl;
  wire mux_354_nl;
  wire or_717_nl;
  wire or_710_nl;
  wire mux_361_nl;
  wire nor_581_nl;
  wire nor_582_nl;
  wire mux_364_nl;
  wire mux_363_nl;
  wire or_740_nl;
  wire or_739_nl;
  wire or_738_nl;
  wire or_742_nl;
  wire nand_19_nl;
  wire mux_372_nl;
  wire mux_371_nl;
  wire or_752_nl;
  wire or_751_nl;
  wire or_750_nl;
  wire mux_375_nl;
  wire nand_20_nl;
  wire mux_386_nl;
  wire mux_385_nl;
  wire mux_384_nl;
  wire mux_383_nl;
  wire mux_382_nl;
  wire mux_381_nl;
  wire mux_380_nl;
  wire mux_379_nl;
  wire mux_378_nl;
  wire mux_377_nl;
  wire mux_376_nl;
  wire or_753_nl;
  wire mux_374_nl;
  wire or_743_nl;
  wire nor_586_nl;
  wire mux_395_nl;
  wire or_772_nl;
  wire mux_394_nl;
  wire mux_393_nl;
  wire or_771_nl;
  wire or_770_nl;
  wire nor_587_nl;
  wire mux_392_nl;
  wire or_764_nl;
  wire mux_391_nl;
  wire mux_390_nl;
  wire or_763_nl;
  wire mux_389_nl;
  wire mux_388_nl;
  wire or_762_nl;
  wire or_761_nl;
  wire or_760_nl;
  wire mux_403_nl;
  wire mux_402_nl;
  wire mux_401_nl;
  wire mux_400_nl;
  wire nor_588_nl;
  wire nor_589_nl;
  wire nor_590_nl;
  wire nor_591_nl;
  wire mux_399_nl;
  wire mux_398_nl;
  wire mux_397_nl;
  wire nor_592_nl;
  wire nor_593_nl;
  wire nor_594_nl;
  wire nor_595_nl;
  wire mux_414_nl;
  wire mux_413_nl;
  wire mux_412_nl;
  wire mux_411_nl;
  wire mux_410_nl;
  wire or_810_nl;
  wire mux_409_nl;
  wire mux_408_nl;
  wire or_809_nl;
  wire or_807_nl;
  wire or_805_nl;
  wire nor_385_nl;
  wire mux_431_nl;
  wire mux_430_nl;
  wire mux_429_nl;
  wire nand_24_nl;
  wire mux_428_nl;
  wire mux_427_nl;
  wire nor_386_nl;
  wire mux_426_nl;
  wire mux_425_nl;
  wire mux_424_nl;
  wire nand_23_nl;
  wire nor_387_nl;
  wire mux_423_nl;
  wire mux_422_nl;
  wire mux_421_nl;
  wire nand_22_nl;
  wire and_760_nl;
  wire mux_420_nl;
  wire nor_388_nl;
  wire mux_419_nl;
  wire mux_418_nl;
  wire mux_417_nl;
  wire nand_21_nl;
  wire nor_389_nl;
  wire mux_416_nl;
  wire or_815_nl;
  wire or_812_nl;
  wire or_845_nl;
  wire mux_434_nl;
  wire mux_433_nl;
  wire or_839_nl;
  wire or_835_nl;
  wire or_830_nl;
  wire mux_439_nl;
  wire mux_438_nl;
  wire mux_437_nl;
  wire mux_436_nl;
  wire or_847_nl;
  wire mux_449_nl;
  wire mux_448_nl;
  wire or_855_nl;
  wire mux_447_nl;
  wire or_877_nl;
  wire or_854_nl;
  wire mux_446_nl;
  wire mux_445_nl;
  wire or_853_nl;
  wire mux_444_nl;
  wire or_878_nl;
  wire or_852_nl;
  wire or_851_nl;
  wire mux_443_nl;
  wire or_879_nl;
  wire or_850_nl;
  wire mux_442_nl;
  wire or_849_nl;
  wire mux_441_nl;
  wire or_880_nl;
  wire or_848_nl;
  wire or_881_nl;
  wire or_858_nl;
  wire or_857_nl;
  wire mux_452_nl;
  wire or_862_nl;
  wire or_861_nl;
  wire mux_462_nl;
  wire mux_461_nl;
  wire mux_460_nl;
  wire mux_459_nl;
  wire or_870_nl;
  wire or_869_nl;
  wire or_868_nl;
  wire or_867_nl;
  wire mux_458_nl;
  wire mux_457_nl;
  wire mux_456_nl;
  wire mux_455_nl;
  wire or_865_nl;
  wire or_864_nl;
  wire mux_454_nl;
  wire or_859_nl;
  wire and_576_nl;
  wire and_575_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl;
  wire weight_mem_banks_write_if_for_if_and_35_nl;
  wire weight_mem_banks_write_if_for_if_and_36_nl;
  wire weight_mem_banks_write_if_for_if_and_37_nl;
  wire weight_mem_banks_write_if_for_if_and_38_nl;
  wire weight_mem_banks_write_if_for_if_and_39_nl;
  wire weight_mem_banks_write_if_for_if_and_40_nl;
  wire weight_mem_banks_write_if_for_if_and_41_nl;
  wire weight_mem_banks_write_if_for_if_mux_7_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl;
  wire mux_159_nl;
  wire nor_610_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl;
  wire weight_mem_banks_write_if_for_if_and_28_nl;
  wire weight_mem_banks_write_if_for_if_and_29_nl;
  wire weight_mem_banks_write_if_for_if_and_30_nl;
  wire weight_mem_banks_write_if_for_if_and_31_nl;
  wire weight_mem_banks_write_if_for_if_and_32_nl;
  wire weight_mem_banks_write_if_for_if_and_33_nl;
  wire weight_mem_banks_write_if_for_if_and_34_nl;
  wire weight_mem_banks_write_if_for_if_mux_6_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl;
  wire mux_158_nl;
  wire nor_609_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl;
  wire weight_mem_banks_write_if_for_if_and_21_nl;
  wire weight_mem_banks_write_if_for_if_and_22_nl;
  wire weight_mem_banks_write_if_for_if_and_23_nl;
  wire weight_mem_banks_write_if_for_if_and_24_nl;
  wire weight_mem_banks_write_if_for_if_and_25_nl;
  wire weight_mem_banks_write_if_for_if_and_26_nl;
  wire weight_mem_banks_write_if_for_if_and_27_nl;
  wire weight_mem_banks_write_if_for_if_mux_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl;
  wire mux_157_nl;
  wire nor_608_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl;
  wire weight_mem_banks_write_if_for_if_and_14_nl;
  wire weight_mem_banks_write_if_for_if_and_15_nl;
  wire weight_mem_banks_write_if_for_if_and_16_nl;
  wire weight_mem_banks_write_if_for_if_and_17_nl;
  wire weight_mem_banks_write_if_for_if_and_18_nl;
  wire weight_mem_banks_write_if_for_if_and_19_nl;
  wire weight_mem_banks_write_if_for_if_and_20_nl;
  wire weight_mem_banks_write_if_for_if_mux_4_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl;
  wire mux_156_nl;
  wire nor_607_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl;
  wire weight_mem_banks_write_if_for_if_and_7_nl;
  wire weight_mem_banks_write_if_for_if_and_8_nl;
  wire weight_mem_banks_write_if_for_if_and_9_nl;
  wire weight_mem_banks_write_if_for_if_and_10_nl;
  wire weight_mem_banks_write_if_for_if_and_11_nl;
  wire weight_mem_banks_write_if_for_if_and_12_nl;
  wire weight_mem_banks_write_if_for_if_and_13_nl;
  wire weight_mem_banks_write_if_for_if_mux_3_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl;
  wire mux_155_nl;
  wire nor_606_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl;
  wire weight_mem_banks_write_if_for_if_and_nl;
  wire weight_mem_banks_write_if_for_if_and_1_nl;
  wire weight_mem_banks_write_if_for_if_and_2_nl;
  wire weight_mem_banks_write_if_for_if_and_3_nl;
  wire weight_mem_banks_write_if_for_if_and_4_nl;
  wire weight_mem_banks_write_if_for_if_and_5_nl;
  wire weight_mem_banks_write_if_for_if_and_6_nl;
  wire weight_mem_banks_write_if_for_if_mux_2_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl;
  wire mux_154_nl;
  wire nor_605_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_1_nl;
  wire weight_mem_banks_write_if_for_if_mux_54_nl;
  wire mux_153_nl;
  wire nor_604_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_nl;
  wire weight_mem_banks_write_if_for_if_mux_53_nl;
  wire mux_152_nl;
  wire nor_603_nl;
  wire rva_out_reg_data_mux_36_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_21_nl;
  wire rva_out_reg_data_mux_37_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_22_nl;
  wire rva_out_reg_data_mux_38_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_23_nl;
  wire PECore_PushAxiRsp_if_else_mux_27_nl;
  wire rva_out_reg_data_mux_40_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_24_nl;
  wire PECore_PushAxiRsp_if_else_mux_28_nl;
  wire rva_out_reg_data_mux_39_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl;
  wire mux_568_nl;
  wire mux_567_nl;
  wire mux_566_nl;
  wire[3:0] mux1h_nl;
  wire not_2446_nl;
  wire[3:0] mux1h_8_nl;
  wire not_2368_nl;
  wire[1:0] mux1h_9_nl;
  wire not_2448_nl;
  wire[3:0] mux1h_10_nl;
  wire not_2370_nl;
  wire mux1h_2_nl;
  wire[6:0] mux1h_11_nl;
  wire not_2449_nl;
  wire mux_32_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_61_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_86_nl;
  wire not_2357_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_66_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_87_nl;
  wire not_2359_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_71_nl;
  wire not_2360_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_88_nl;
  wire not_2361_nl;
  wire mux_34_nl;
  wire or_211_nl;
  wire[1:0] weight_mem_banks_load_store_for_else_mux1h_76_nl;
  wire not_2362_nl;
  wire[5:0] weight_mem_banks_load_store_for_else_mux1h_89_nl;
  wire not_2363_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_80_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_90_nl;
  wire not_2365_nl;
  wire mux_38_nl;
  wire nor_494_nl;
  wire mux_37_nl;
  wire nor_495_nl;
  wire mux_36_nl;
  wire mux_35_nl;
  wire nor_496_nl;
  wire mux_493_nl;
  wire weight_mem_banks_load_store_for_else_or_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_85_nl;
  wire[6:0] mux_494_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_or_1_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_91_nl;
  wire and_687_nl;
  wire not_2367_nl;
  wire mux1h_5_nl;
  wire[6:0] mux1h_12_nl;
  wire not_2450_nl;
  wire mux1h_6_nl;
  wire[6:0] mux1h_13_nl;
  wire not_2451_nl;
  wire mux1h_7_nl;
  wire[6:0] mux1h_14_nl;
  wire not_2452_nl;
  wire mux_5_nl;
  wire mux_593_nl;
  wire mux_592_nl;
  wire nor_743_nl;
  wire mux_591_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_130_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_237_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_128_nl;
  wire[1:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_135_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_265_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_136_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl;
  wire mux_607_nl;
  wire mux_606_nl;
  wire nor_745_nl;
  wire mux_605_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_129_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_267_nl;
  wire mux_614_nl;
  wire mux_613_nl;
  wire nor_746_nl;
  wire mux_612_nl;
  wire mux_617_nl;
  wire or_1188_nl;
  wire or_1186_nl;
  wire mux_616_nl;
  wire mux_615_nl;
  wire or_1185_nl;
  wire or_1184_nl;
  wire or_1183_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_107_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_123_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_106_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_122_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_133_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_275_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_134_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_276_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_138_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_278_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_137_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_277_nl;
  wire[3:0] while_if_while_if_and_27_nl;
  wire[3:0] while_if_while_if_and_35_nl;
  wire[3:0] while_if_while_if_and_37_nl;
  wire[6:0] while_if_while_if_and_33_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_110_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_126_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_145_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_281_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_146_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_282_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_109_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_125_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_147_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_283_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_148_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_284_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_108_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_279_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_124_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_280_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_139_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_147_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_140_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_162_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_18_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_mux_25_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_mux_26_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_27_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_20_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_28_nl;
  wire mux1h_1_nl;
  wire mux1h_15_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_131_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_132_nl;
  wire[1:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_141_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl;
  wire[1:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_142_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_273_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_143_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_271_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_144_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_274_nl;
  wire[6:0] while_if_while_if_and_39_nl;
  wire[6:0] while_if_while_if_and_38_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_19_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_30_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_29_nl;
  wire mux_564_nl;
  wire mux_563_nl;
  wire or_1125_nl;
  wire or_1124_nl;
  wire or_1123_nl;
  wire mux_576_nl;
  wire mux_575_nl;
  wire or_1141_nl;
  wire or_1140_nl;
  wire or_1139_nl;
  wire or_1144_nl;
  wire mux_589_nl;
  wire and_1642_nl;
  wire mux_588_nl;
  wire mux_587_nl;
  wire and_1643_nl;
  wire and_1644_nl;
  wire and_1645_nl;
  wire mux_603_nl;
  wire and_1652_nl;
  wire mux_602_nl;
  wire mux_601_nl;
  wire and_1653_nl;
  wire and_1654_nl;
  wire and_1655_nl;
  wire mux_610_nl;
  wire and_1657_nl;
  wire mux_609_nl;
  wire mux_608_nl;
  wire and_1658_nl;
  wire and_1659_nl;
  wire and_1660_nl;
  wire mux_550_nl;
  wire or_1048_nl;
  wire nor_638_nl;
  wire mux_580_nl;
  wire mux_579_nl;
  wire mux_578_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (~ reg_rva_in_reg_rw_sva_2_cse);
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0];
  wire  nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a = PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2
      & reg_rva_in_reg_rw_sva_2_cse;
  wire [2:0] nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s = weight_write_addrs_lpi_1_dfm_1_2[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s = {(weight_read_addrs_6_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_4[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s = weight_read_addrs_7_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s = {(weight_read_addrs_2_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s = {(weight_read_addrs_4_14_2_lpi_1_dfm_1_1[0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[1:0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s = weight_read_addrs_3_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s = weight_read_addrs_5_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s = weight_read_addrs_1_lpi_1_dfm_1_1[2:0];
  wire [255:0] nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff;
  assign nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff
      = {15'b000000000000000 , act_port_reg_data_240_224_sva_dfm_1_2 , 15'b000000000000000
      , act_port_reg_data_208_192_sva_dfm_1_2 , 15'b000000000000000 , act_port_reg_data_176_160_sva_dfm_1_2
      , 15'b000000000000000 , act_port_reg_data_144_128_sva_dfm_1_1 , 15'b000000000000000
      , act_port_reg_data_112_96_sva_dfm_1_1 , 15'b000000000000000 , act_port_reg_data_80_64_sva_dfm_1_1
      , 15'b000000000000000 , act_port_reg_data_48_32_sva_dfm_1_1 , 15'b000000000000000
      , act_port_reg_data_16_0_sva_dfm_1_2};
  wire weight_port_read_out_data_mux_4_nl;
  wire weight_port_read_out_data_mux_149_nl;
  wire weight_port_read_out_data_mux_2_nl;
  wire weight_port_read_out_data_mux_148_nl;
  wire weight_port_read_out_data_mux_nl;
  wire weight_port_read_out_data_mux_147_nl;
  wire [127:0] nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign weight_port_read_out_data_mux_149_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_26_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign weight_port_read_out_data_mux_4_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2,
      weight_port_read_out_data_mux_149_nl, fsm_output);
  assign weight_port_read_out_data_mux_148_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_25_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign weight_port_read_out_data_mux_2_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2,
      weight_port_read_out_data_mux_148_nl, fsm_output);
  assign weight_port_read_out_data_mux_147_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_24_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign weight_port_read_out_data_mux_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2,
      weight_port_read_out_data_mux_147_nl, fsm_output);
  assign nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun
      = {rva_out_reg_data_127_120_sva_dfm_4_5 , rva_out_reg_data_119_112_sva_dfm_4_5_rsp_0
      , rva_out_reg_data_119_112_sva_dfm_4_5_rsp_1 , rva_out_reg_data_111_104_sva_dfm_4_5_rsp_0
      , rva_out_reg_data_111_104_sva_dfm_4_5_rsp_1 , rva_out_reg_data_103_96_sva_dfm_4_5_7_4
      , rva_out_reg_data_103_96_sva_dfm_4_5_3_0 , rva_out_reg_data_95_88_sva_dfm_4_5_rsp_0
      , rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_0 , rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_1
      , rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_2 , rva_out_reg_data_87_80_sva_dfm_4_5_rsp_0
      , rva_out_reg_data_87_80_sva_dfm_4_5_rsp_1 , rva_out_reg_data_79_72_sva_dfm_4_5
      , rva_out_reg_data_71_64_sva_dfm_4_5 , rva_out_reg_data_63_sva_dfm_4_5 , rva_out_reg_data_62_56_sva_dfm_4_5
      , rva_out_reg_data_55_48_sva_dfm_4_5 , rva_out_reg_data_47_sva_dfm_4_5 , rva_out_reg_data_46_40_sva_dfm_4_5
      , rva_out_reg_data_39_36_sva_dfm_4_5_3 , rva_out_reg_data_39_36_sva_dfm_4_5_2_0
      , rva_out_reg_data_35_32_sva_dfm_4_5 , PECore_PushAxiRsp_if_mux1h_17 , PECore_PushAxiRsp_if_mux1h_16_5_3
      , PECore_PushAxiRsp_if_mux1h_16_2_0 , PECore_PushAxiRsp_if_mux1h_15 , PECore_PushAxiRsp_if_mux1h_14_6
      , PECore_PushAxiRsp_if_mux1h_14_5 , PECore_PushAxiRsp_if_mux1h_14_4_3 , PECore_PushAxiRsp_if_mux1h_14_2_0
      , weight_port_read_out_data_mux_4_nl , PECore_PushAxiRsp_if_mux1h_12_6 , PECore_PushAxiRsp_if_mux1h_12_5_0
      , weight_port_read_out_data_mux_2_nl , PECore_PushAxiRsp_if_mux1h_10_6 , PECore_PushAxiRsp_if_mux1h_10_5_0
      , weight_port_read_out_data_mux_nl};
  PECore_mgc_muladd1 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_cst(32'sd1),
  .signd_cst(32'sd0),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd11),
  .add_axb(32'sd1),
  .add_c(32'sd1),
  .add_d(32'sd1),
  .use_const(32'sd1)) PEManager_15U_GetWeightAddr_else_acc_4_cmp (
      .a(pe_config_output_counter_sva),
      .b(pe_manager_num_input_sva),
      .c(pe_config_input_counter_sva),
      .cst(1'b0),
      .z(PEManager_15U_GetWeightAddr_else_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_for_1_lshift_rg (
      .a(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a),
      .s(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_write_arbxbar_xbar_for_lshift_rg (
      .a(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a),
      .s(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s[2:0]),
      .z(weight_mem_write_arbxbar_xbar_for_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi PECore_PECoreRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(fsm_output)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi PECore_PECoreRun_input_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_oswt_pff(and_570_rmff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi PECore_PECoreRun_act_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(reg_act_port_Push_mioi_iswt0_cse),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff(nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[255:0]),
      .act_port_Push_mioi_oswt_pff(and_572_rmff)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi PECore_PECoreRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_oswt_pff(and_570_rmff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi PECore_PECoreRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun[127:0]),
      .rva_out_Push_mioi_oswt_pff(and_568_cse)
    );
  PECore_PECore_PECoreRun_wait_dp PECore_PECoreRun_wait_dp_inst (
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .PECoreRun_wen(PECoreRun_wen),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg(and_566_rmff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg(and_563_rmff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg(and_558_rmff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg(and_554_rmff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg(and_549_rmff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg(and_545_rmff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg(and_541_rmff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg(and_537_rmff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_cgo(reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_56_cse),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg(and_533_rmff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_1(reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_63_cse),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg_1(and_530_rmff)
    );
  PECore_PECore_PECoreRun_staller PECore_PECoreRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp)
    );
  PECore_PECore_PECoreRun_PECoreRun_fsm PECore_PECoreRun_PECoreRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .fsm_output(fsm_output)
    );
  assign weight_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_96);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign weight_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_96);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign weight_mem_banks_read_1_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_98);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign weight_mem_banks_read_1_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_98);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign weight_mem_banks_read_1_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_100);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 );
  assign weight_mem_banks_read_1_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_100);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign weight_mem_banks_read_1_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_102);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 );
  assign weight_mem_banks_read_1_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_102);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign weight_mem_banks_read_1_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_104);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 );
  assign weight_mem_banks_read_1_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_104);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign weight_mem_banks_read_1_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_106);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 );
  assign weight_mem_banks_read_1_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_106);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign weight_mem_banks_read_1_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_92);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 );
  assign weight_mem_banks_read_1_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_92);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign weight_mem_banks_read_1_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_94);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 );
  assign weight_mem_banks_read_1_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_94);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign weight_mem_banks_write_if_for_if_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_189);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 );
  assign weight_mem_banks_write_if_for_if_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_189);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign weight_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_190);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 );
  assign weight_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_190);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign weight_mem_banks_write_if_for_if_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_192);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 );
  assign weight_mem_banks_write_if_for_if_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_192);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1
      = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1
      = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign weight_mem_banks_read_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_193);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 );
  assign weight_mem_banks_read_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_193);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign weight_mem_banks_write_if_for_if_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_195);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 );
  assign weight_mem_banks_write_if_for_if_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_195);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2
      = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2
      = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign weight_mem_banks_read_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_196);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 );
  assign weight_mem_banks_read_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_196);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign weight_mem_banks_write_if_for_if_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_198);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 );
  assign weight_mem_banks_write_if_for_if_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_198);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3
      = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3
      = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign weight_mem_banks_read_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_199);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 );
  assign weight_mem_banks_read_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_199);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign weight_mem_banks_write_if_for_if_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_200);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 );
  assign weight_mem_banks_write_if_for_if_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_200);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4
      = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4
      = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign weight_mem_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_201);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 );
  assign weight_mem_banks_read_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_201);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign weight_mem_banks_write_if_for_if_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_202);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 );
  assign weight_mem_banks_write_if_for_if_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_202);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5
      = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5
      = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign weight_mem_banks_read_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_203);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 );
  assign weight_mem_banks_read_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_203);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign weight_mem_banks_write_if_for_if_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_205);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 );
  assign weight_mem_banks_write_if_for_if_mux_33_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_205);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6
      = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6
      = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign weight_mem_banks_read_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_206);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 );
  assign weight_mem_banks_read_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_206);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign weight_mem_banks_write_if_for_if_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_208);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 );
  assign weight_mem_banks_write_if_for_if_mux_37_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_208);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7
      = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7
      = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign weight_mem_banks_read_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_209);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 );
  assign weight_mem_banks_read_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_209);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign input_mem_banks_write_1_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_219);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 );
  assign input_mem_banks_write_1_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_219);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8
      = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_3 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8
      = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign input_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_216);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 );
  assign input_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_216);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign input_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_228);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 );
  assign input_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_228);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9
      = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_1 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9
      = input_mem_banks_write_if_for_if_mux_1_cse;
  assign input_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_230);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 );
  assign input_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_230);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign and_527_cse = and_dcpl_33 & PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  assign and_530_rmff = (and_dcpl_528 | and_527_cse | and_dcpl_524) & fsm_output;
  assign and_533_rmff = (and_dcpl_528 | (while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_8) | and_dcpl_524) & fsm_output;
  assign or_334_nl = (weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & while_stage_0_7) | and_tmp_1;
  assign or_333_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3)
      | (~ while_stage_0_7))) | and_tmp_1;
  assign mux_112_nl = MUX_s_1_2_2(or_334_nl, or_333_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_537_rmff = (mux_112_nl | and_dcpl_534) & fsm_output;
  assign or_338_nl = (weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & while_stage_0_7) | and_tmp_2;
  assign or_337_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3)
      | (~ while_stage_0_7))) | and_tmp_2;
  assign mux_114_nl = MUX_s_1_2_2(or_338_nl, or_337_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_541_rmff = (mux_114_nl | and_dcpl_537) & fsm_output;
  assign or_343_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_3;
  assign or_342_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2)))
      | and_tmp_3;
  assign mux_117_nl = MUX_s_1_2_2(or_343_nl, or_342_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_118_nl = MUX_s_1_2_2(and_tmp_3, mux_117_nl, while_stage_0_6);
  assign and_545_rmff = (mux_118_nl | and_dcpl_202) & fsm_output;
  assign or_350_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_5;
  assign or_882_nl = (~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1)) | and_tmp_5;
  assign mux_121_nl = MUX_s_1_2_2(or_350_nl, or_882_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_122_nl = MUX_s_1_2_2(and_tmp_5, mux_121_nl, while_stage_0_6);
  assign and_549_rmff = (mux_122_nl | and_dcpl_200) & fsm_output;
  assign or_356_nl = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_7;
  assign or_355_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse)))
      | and_tmp_7;
  assign mux_124_nl = MUX_s_1_2_2(or_356_nl, or_355_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_125_nl = MUX_s_1_2_2(and_tmp_7, mux_124_nl, while_stage_0_6);
  assign and_554_rmff = (mux_125_nl | and_dcpl_545) & fsm_output;
  assign or_361_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_8;
  assign or_883_nl = (~((~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1)) | and_tmp_8;
  assign mux_128_nl = MUX_s_1_2_2(or_361_nl, or_883_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_129_nl = MUX_s_1_2_2(and_tmp_8, mux_128_nl, while_stage_0_6);
  assign and_558_rmff = (mux_129_nl | and_dcpl_195) & fsm_output;
  assign or_367_nl = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | mux_tmp_132;
  assign or_366_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse)))
      | mux_tmp_132;
  assign mux_133_nl = MUX_s_1_2_2(or_367_nl, or_366_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_134_nl = MUX_s_1_2_2(mux_tmp_132, mux_133_nl, while_stage_0_6);
  assign and_563_rmff = (mux_134_nl | and_dcpl_192) & fsm_output;
  assign or_373_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_11;
  assign or_884_nl = (~((~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1)) | and_tmp_11;
  assign mux_136_nl = MUX_s_1_2_2(or_373_nl, or_884_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_137_nl = MUX_s_1_2_2(and_tmp_11, mux_136_nl, while_stage_0_6);
  assign and_566_rmff = (mux_137_nl | and_dcpl_189) & fsm_output;
  assign and_1209_itm = PECore_UpdateFSM_switch_lp_nor_7_itm_1 & PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      & pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign and_809_itm = pe_config_is_zero_first_sva & PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      & pe_manager_zero_active_sva;
  assign and_1089_cse = PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign mux_654_nl = MUX_s_1_2_2(and_1209_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_809_itm);
  assign and_1088_nl = start_PopNB_mioi_data_rsc_z_mxwt & start_PopNB_mioi_return_rsc_z_mxwt
      & PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign mux_146_nl = MUX_s_1_2_2(mux_654_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_1088_nl);
  assign mux_495_nl = MUX_s_1_2_2(and_1209_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_809_itm);
  assign mux_142_nl = MUX_s_1_2_2(mux_495_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_1089_cse);
  assign mux_147_nl = MUX_s_1_2_2(mux_146_nl, mux_142_nl, or_380_cse);
  assign mux_663_nl = MUX_s_1_2_2(and_1209_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_809_itm);
  assign mux_662_nl = MUX_s_1_2_2(mux_663_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_1089_cse);
  assign or_378_nl = pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]);
  assign mux_143_nl = MUX_s_1_2_2(mux_662_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_378_nl);
  assign or_377_nl = (state_2_1_sva!=2'b10) | state_0_sva;
  assign mux_144_nl = MUX_s_1_2_2(mux_143_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_377_nl);
  assign mux_145_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_nor_7_itm_1, mux_144_nl,
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign mux_148_nl = MUX_s_1_2_2(mux_147_nl, mux_145_nl, PECore_UpdateFSM_switch_lp_equal_tmp_5_1);
  assign mux_149_nl = MUX_s_1_2_2(mux_148_nl, state_0_sva, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_150_nl = MUX_s_1_2_2(or_380_cse, mux_149_nl, while_stage_0_3);
  assign or_376_nl = while_stage_0_3 | (state_2_1_sva!=2'b00) | state_0_sva;
  assign or_375_nl = (state_2_1_sva_dfm_1!=2'b00);
  assign mux_151_nl = MUX_s_1_2_2(mux_150_nl, or_376_nl, or_375_nl);
  assign and_570_rmff = (~ mux_151_nl) & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign and_572_rmff = while_stage_0_12 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10)
      & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10;
  assign PECore_DecodeAxiRead_switch_lp_and_2_cse = PECoreRun_wen & and_dcpl_5 &
      and_dcpl_2 & (~ input_read_req_valid_lpi_1_dfm_1_9);
  assign rva_out_reg_data_and_22_cse = PECoreRun_wen & and_dcpl_5 & and_dcpl_2 &
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 | rva_in_reg_rw_sva_st_9)) &
      (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_9 | input_read_req_valid_lpi_1_dfm_1_9));
  assign rva_out_reg_data_and_147_enex5 = rva_out_reg_data_and_22_cse & reg_rva_out_reg_data_15_9_sva_dfm_9_enexo;
  assign rva_out_reg_data_and_148_enex5 = rva_out_reg_data_and_22_cse & reg_rva_out_reg_data_23_17_sva_dfm_7_enexo;
  assign rva_out_reg_data_and_149_enex5 = rva_out_reg_data_and_22_cse & reg_rva_out_reg_data_30_25_sva_dfm_7_enexo;
  assign rva_out_reg_data_and_25_cse = PECoreRun_wen & and_dcpl_5;
  assign rva_out_reg_data_and_150_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_127_120_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_151_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_79_72_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_152_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_71_64_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_153_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_154_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_155_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_156_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo;
  assign input_mem_banks_read_read_data_and_cse = PECoreRun_wen & and_dcpl_5 & (~
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7) & input_read_req_valid_lpi_1_dfm_1_9;
  assign weight_port_read_out_data_and_123_cse = PECoreRun_wen & and_dcpl_4 & (~
      rva_in_reg_rw_sva_st_1_9) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
  assign rva_out_reg_data_and_cse = PECoreRun_wen & (~((~(while_stage_0_12 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10))
      | rva_in_reg_rw_sva_10 | (~ fsm_output)));
  assign input_mem_banks_read_read_data_and_47_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo;
  assign input_mem_banks_read_read_data_and_48_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo;
  assign input_mem_banks_read_read_data_and_49_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo;
  assign input_mem_banks_read_read_data_and_50_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo;
  assign rva_in_reg_rw_and_cse = PECoreRun_wen & while_stage_0_11;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_cse = PECoreRun_wen & and_dcpl_4
      & (~(rva_in_reg_rw_sva_st_1_9 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7))
      & (~ rva_in_reg_rw_sva_9) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 &
      (~ input_read_req_valid_lpi_1_dfm_1_9);
  assign act_port_reg_data_and_cse = PECoreRun_wen & and_dcpl_24 & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  assign act_port_reg_data_and_19_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_16_0_sva_dfm_1_1_enexo;
  assign act_port_reg_data_and_20_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_240_224_sva_dfm_1_1_enexo;
  assign and_1224_cse = (PECore_UpdateFSM_switch_lp_equal_tmp_2_10 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
      | (~ while_stage_0_12) | ((~ PECore_RunMac_PECore_RunMac_if_and_svs_st_9) &
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9)) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)
      & PECoreRun_wen & while_stage_0_11 & (PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9
      | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9));
  assign act_port_reg_data_and_21_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_208_192_sva_dfm_1_1_enexo;
  assign act_port_reg_data_and_22_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_176_160_sva_dfm_1_1_enexo;
  assign PECore_PushOutput_if_and_cse = PECoreRun_wen & and_dcpl_24;
  assign PECore_RunMac_if_and_cse = PECoreRun_wen & and_1462_cse;
  assign while_if_and_6_cse = PECoreRun_wen & while_stage_0_10;
  assign rva_in_reg_rw_and_2_cse = PECoreRun_wen & and_dcpl_29;
  assign PECore_RunMac_if_and_1_cse = PECoreRun_wen & (and_dcpl_30 | and_dcpl_346);
  assign while_if_and_7_cse = PECoreRun_wen & while_stage_0_9;
  assign PECore_RunMac_if_and_2_cse = PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
      & rva_in_reg_rw_sva_st_1_6)) & while_stage_0_8;
  assign while_if_and_8_cse = PECoreRun_wen & while_stage_0_8;
  assign input_mem_banks_read_1_read_data_and_enex5 = PECoreRun_wen & and_527_cse
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  assign mux_1_nl = MUX_s_1_2_2(mux_tmp, (~ weight_mem_run_3_for_land_2_lpi_1_dfm_2),
      while_stage_0_7);
  assign or_6_nl = while_stage_0_7 | mux_tmp;
  assign mux_2_nl = MUX_s_1_2_2(mux_1_nl, or_6_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign weight_port_read_out_data_and_enex5 = PECoreRun_wen & (~(or_dcpl_221 | (~
      weight_mem_run_3_for_land_2_lpi_1_dfm_3) | (~ fsm_output))) & mux_2_nl & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  assign weight_mem_run_3_for_aelse_and_cse = PECoreRun_wen & while_stage_0_7;
  assign weight_port_read_out_data_and_1_cse = PECoreRun_wen & (~(or_dcpl_221 | (~
      weight_mem_run_3_for_land_3_lpi_1_dfm_3)));
  assign weight_port_read_out_data_and_190_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  assign data_in_tmp_operator_2_for_and_1_cse = PECoreRun_wen & and_dcpl_33 & weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  assign weight_port_read_out_data_and_191_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001;
  assign weight_port_read_out_data_and_192_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002;
  assign weight_port_read_out_data_and_193_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003;
  assign weight_port_read_out_data_and_194_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004;
  assign weight_port_read_out_data_and_195_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005;
  assign weight_port_read_out_data_and_196_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006;
  assign weight_port_read_out_data_and_197_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007;
  assign weight_port_read_out_data_and_198_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008;
  assign weight_port_read_out_data_and_199_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009;
  assign weight_port_read_out_data_and_200_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010;
  assign weight_port_read_out_data_and_201_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011;
  assign weight_port_read_out_data_and_202_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012;
  assign weight_port_read_out_data_and_203_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013;
  assign weight_port_read_out_data_and_204_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014;
  assign weight_port_read_out_data_and_16_cse = PECoreRun_wen & (~(or_dcpl_221 |
      (~ weight_mem_run_3_for_land_5_lpi_1_dfm_3)));
  assign weight_port_read_out_data_and_205_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  assign data_in_tmp_operator_2_for_and_16_cse = PECoreRun_wen & and_dcpl_33 & weight_mem_run_3_for_land_5_lpi_1_dfm_2;
  assign weight_port_read_out_data_and_206_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001;
  assign weight_port_read_out_data_and_207_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002;
  assign weight_port_read_out_data_and_208_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003;
  assign weight_port_read_out_data_and_209_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004;
  assign weight_port_read_out_data_and_210_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005;
  assign weight_port_read_out_data_and_211_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006;
  assign weight_port_read_out_data_and_212_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007;
  assign weight_port_read_out_data_and_213_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008;
  assign weight_port_read_out_data_and_214_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009;
  assign weight_port_read_out_data_and_215_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010;
  assign weight_port_read_out_data_and_216_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011;
  assign weight_port_read_out_data_and_217_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012;
  assign weight_port_read_out_data_and_218_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013;
  assign weight_port_read_out_data_and_219_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014;
  assign weight_port_read_out_data_and_31_enex5 = PECoreRun_wen & (~(or_dcpl_221
      | (~ weight_mem_run_3_for_land_4_lpi_1_dfm_3) | (~ fsm_output))) & ((~ while_stage_0_7)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)) & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000;
  assign PECore_RunMac_if_and_3_cse = PECoreRun_wen & nand_32_cse & while_stage_0_7;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2:1]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      | (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1:0]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_or_1_cse = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3) | ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_1147_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_dcpl);
  assign and_1148_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_1_cse & (~
      or_dcpl);
  assign and_1149_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      & (~ or_dcpl);
  assign and_1150_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1
      & (~ or_dcpl);
  assign and_1151_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      & (~ or_dcpl);
  assign and_1152_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      & (~ or_dcpl);
  assign nor_626_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl);
  assign and_1156_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_1_cse & (~
      or_dcpl_296);
  assign and_1157_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      & (~ or_dcpl_296);
  assign and_1158_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      & (~ or_dcpl_296);
  assign and_1159_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      & (~ or_dcpl_296);
  assign and_1160_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      & (~ or_dcpl_296);
  assign nor_627_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl_296);
  assign rva_in_reg_rw_and_3_cse = PECoreRun_wen & and_dcpl_48;
  assign weight_mem_banks_read_1_read_data_and_8_cse = PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign input_mem_banks_read_1_read_data_and_1_enex5 = PECoreRun_wen & reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  assign weight_port_read_out_data_and_136_cse = PECoreRun_wen & ((weight_mem_run_3_for_land_1_lpi_1_dfm_3
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5))
      | while_and_40_tmp) & while_stage_0_7 & fsm_output & (~(mux_6_itm & while_stage_0_6));
  assign weight_mem_run_3_for_aelse_and_4_cse = PECoreRun_wen & while_stage_0_6;
  assign weight_port_read_out_data_and_41_cse = PECoreRun_wen & weight_mem_run_3_for_land_7_lpi_1_dfm_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7;
  assign weight_port_read_out_data_and_145_cse = PECoreRun_wen & (~((~(weight_mem_run_3_for_land_2_lpi_1_dfm_2
      & while_stage_0_7)) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ fsm_output))) & mux_tmp;
  assign or_18_nl = (~ weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp) | (~
      while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_8_nl = MUX_s_1_2_2(or_18_nl, or_tmp_7, while_stage_0_6);
  assign weight_port_read_out_data_and_159_cse = PECoreRun_wen & (~(or_dcpl_231 |
      (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2) | (~ fsm_output))) & mux_8_nl;
  assign weight_port_read_out_data_and_85_cse = PECoreRun_wen & (~ or_dcpl_233);
  assign weight_port_read_out_data_7_15_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), weight_port_read_out_data_7_15_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_143_itm_2 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign xor_1_cse = (weight_read_addrs_7_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[2]);
  assign and_1244_cse = (xor_1_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_port_read_out_data_7_14_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), weight_port_read_out_data_7_14_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign nor_681_cse = ~((weight_read_addrs_7_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_516_nl = MUX_s_1_2_2((weight_read_addrs_7_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_7_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_7_lpi_1_dfm_3_2_0[0]);
  assign mux_517_cse = MUX_s_1_2_2(mux_516_nl, nor_681_cse, weight_read_addrs_7_lpi_1_dfm_3_2_0[2]);
  assign and_1249_cse = (mux_517_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_port_read_out_data_7_13_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), weight_port_read_out_data_7_13_sva_dfm_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign and_1254_cse = (xor_1_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_port_read_out_data_7_12_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]), weight_port_read_out_data_7_12_sva_dfm_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_11_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]), weight_port_read_out_data_7_11_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_143_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_10_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]), weight_port_read_out_data_7_10_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_100_itm_1 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_9_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]), weight_port_read_out_data_7_9_sva_dfm_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign and_1274_cse = (mux_517_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_port_read_out_data_7_8_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]), weight_port_read_out_data_7_8_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_143_itm_2 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign and_1280_cse = (and_1244_cse | weight_mem_run_3_for_5_and_143_itm_2 | weight_mem_run_3_for_5_and_134_itm_2
      | weight_mem_run_3_for_5_and_140_itm_2) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & weight_mem_run_3_for_aelse_and_cse;
  assign weight_port_read_out_data_7_7_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]), weight_port_read_out_data_7_7_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_143_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign and_1285_cse = (and_1249_cse | or_dcpl_337 | or_dcpl_323) & fsm_output &
      (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & weight_mem_run_3_for_aelse_and_cse;
  assign weight_port_read_out_data_7_6_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]), weight_port_read_out_data_7_6_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_143_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_5_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]), weight_port_read_out_data_7_5_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_143_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_4_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]), weight_port_read_out_data_7_4_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_143_itm_2 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_3_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]), weight_port_read_out_data_7_3_sva_dfm_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_100_itm_1 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_2_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]), weight_port_read_out_data_7_2_sva_dfm_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_100_itm_1 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_143_itm_2 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_1_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]), weight_port_read_out_data_7_1_sva_dfm_1,
      {weight_mem_run_3_for_5_and_156 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_134_itm_2
      , weight_mem_run_3_for_5_and_143_itm_2 , weight_mem_run_3_for_5_asn_453 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_0_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]),
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9, weight_port_read_out_data_7_0_sva_dfm_1,
      {weight_mem_run_3_for_5_and_152 , weight_mem_run_3_for_5_asn_447 , weight_mem_run_3_for_5_asn_449
      , weight_mem_run_3_for_5_and_100_itm_1 , weight_mem_run_3_for_5_asn_451 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_135_itm_1 , weight_mem_run_3_for_5_and_136_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_15_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), weight_port_read_out_data_5_15_sva_dfm_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , weight_mem_run_3_for_5_and_12_itm_1 , weight_mem_run_3_for_5_asn_459
      , reg_weight_mem_run_3_for_5_and_14_itm_1_cse , reg_weight_mem_run_3_for_5_and_15_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_16_itm_1_cse , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign nor_690_cse = ~((weight_read_addrs_5_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_534_nl = MUX_s_1_2_2((weight_read_addrs_5_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_5_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_5_lpi_1_dfm_3_2_0[0]);
  assign mux_535_nl = MUX_s_1_2_2(mux_534_nl, nor_690_cse, weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign and_1324_cse = (mux_535_nl | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_port_read_out_data_5_14_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), weight_port_read_out_data_5_14_sva_dfm_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , weight_mem_run_3_for_5_and_7_itm_1 , reg_weight_mem_run_3_for_5_and_16_itm_1_cse
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_372_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_6_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_380_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_384_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_4_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_389_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_390_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_2_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_cse = PECoreRun_wen
      & not_tmp_29 & while_stage_0_6;
  assign and_797_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  assign and_798_cse = weight_mem_read_arbxbar_arbiters_next_7_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign and_799_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  assign and_800_cse = weight_mem_read_arbxbar_arbiters_next_6_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign weight_read_addrs_and_5_cse = PECoreRun_wen & (((~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]))
      & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1)
      | (weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
      & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7])))) & and_dcpl_83;
  assign weight_read_addrs_and_28_enex5 = weight_read_addrs_and_5_cse & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse = PECoreRun_wen & and_dcpl_92;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse
      & (reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_enexo | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1);
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse = PECoreRun_wen & and_dcpl_94;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse
      & (reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_enexo_1 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2_enexo
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo_1
      | reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo);
  assign while_if_and_11_cse = PECoreRun_wen & while_stage_0_5;
  assign weight_mem_read_arbxbar_arbiters_next_and_cse = PECoreRun_wen & fsm_output;
  assign weight_mem_read_arbxbar_arbiters_next_and_49_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_113_cse | or_dcpl_75);
  assign weight_mem_read_arbxbar_arbiters_next_and_55_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_120_cse | or_dcpl_75);
  assign weight_mem_read_arbxbar_arbiters_next_and_61_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_127_cse | or_dcpl_75);
  assign weight_mem_read_arbxbar_arbiters_next_and_67_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_134_cse | or_dcpl_75);
  assign weight_mem_read_arbxbar_arbiters_next_and_73_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & or_dcpl_80;
  assign weight_mem_read_arbxbar_arbiters_next_and_78_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_148_cse | or_dcpl_75);
  assign weight_mem_read_arbxbar_arbiters_next_and_84_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (((~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])))
      & nor_427_cse & nor_428_cse) | or_dcpl_75);
  assign weight_mem_read_arbxbar_arbiters_next_and_90_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_162_cse | or_dcpl_75);
  assign weight_read_addrs_and_7_cse = PECoreRun_wen & (and_dcpl_170 | and_dcpl_169
      | and_dcpl_168 | and_dcpl_167 | and_dcpl_166 | and_dcpl_165 | and_dcpl_164
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | and_dcpl_163) & while_stage_0_4;
  assign weight_write_data_data_and_cse = PECoreRun_wen & ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7:6]!=2'b00))
      & and_dcpl_172;
  assign weight_write_data_data_and_48_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_49_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_50_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_51_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_52_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_53_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_54_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_55_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_56_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_57_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_58_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_59_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_60_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_61_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_62_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_63_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_addrs_and_enex5 = weight_write_data_data_and_cse & reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  assign weight_mem_write_arbxbar_xbar_for_1_for_and_cse = PECoreRun_wen & and_dcpl_172;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
      = PECoreRun_wen & and_dcpl_180;
  assign PECore_RunFSM_switch_lp_and_cse = PECoreRun_wen & while_stage_0_4;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 & and_dcpl_180;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 & and_dcpl_180;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12 & and_dcpl_180;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14 & and_dcpl_180;
  assign Arbiter_8U_Roundrobin_pick_1_and_15_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8
      & and_dcpl_180;
  assign Arbiter_8U_Roundrobin_pick_and_cse = PECoreRun_wen & (while_stage_0_4 |
      and_dcpl_600) & fsm_output & or_dcpl_75;
  assign Arbiter_8U_Roundrobin_pick_1_and_22_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9
      & and_dcpl_180;
  assign Arbiter_8U_Roundrobin_pick_1_and_50_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13
      & and_dcpl_180;
  assign Arbiter_8U_Roundrobin_pick_1_and_64_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15
      & and_dcpl_180;
  assign weight_write_data_data_and_16_cse = PECoreRun_wen & and_dcpl_212;
  assign weight_write_data_data_and_64_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_65_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_66_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_67_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_68_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_69_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_70_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_71_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_72_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_73_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_74_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_75_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_76_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_77_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_78_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_79_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  assign weight_write_addrs_and_2_enex5 = weight_write_data_data_and_16_cse & reg_pe_manager_base_input_enexo;
  assign rva_in_reg_rw_and_4_cse = PECoreRun_wen & while_stage_0_3;
  assign weight_read_addrs_and_29_enex5 = weight_write_data_data_and_16_cse & reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  assign state_and_cse = weight_mem_read_arbxbar_arbiters_next_and_cse & nand_88_cse;
  assign and_1341_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & while_stage_0_3;
  assign pe_config_num_manager_and_cse = PECoreRun_wen & (~(or_dcpl_249 | nand_88_cse
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])))));
  assign rva_in_reg_rw_and_5_cse = PECoreRun_wen & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign PECore_UpdateFSM_switch_lp_and_9_cse = PECoreRun_wen & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign pe_config_UpdateManagerCounter_if_if_and_enex5 = PECoreRun_wen & reg_pe_config_num_output_enexo;
  assign PECore_DecodeAxiRead_switch_lp_and_cse = PECoreRun_wen & (~(nand_88_cse
      | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
  assign PECore_DecodeAxiWrite_switch_lp_and_cse = PECoreRun_wen & (~ or_dcpl_256);
  assign and_1374_cse = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
      | (~ while_stage_0_11)) & while_stage_0_12 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10)
      & fsm_output & PECoreRun_wen;
  assign and_1393_cse = ((~(((~(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_8)) & PECore_UpdateFSM_switch_lp_equal_tmp_2_8)
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_8)) | (~ while_stage_0_10) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)
      & PECoreRun_wen & (PECore_UpdateFSM_switch_lp_equal_tmp_2_9 | PECore_RunMac_PECore_RunMac_if_and_svs_st_9)
      & while_stage_0_11;
  assign nor_12_cse = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7));
  assign mux_29_nl = MUX_s_1_2_2(and_1619_cse, mux_tmp_4, nor_12_cse);
  assign weight_mem_banks_load_store_for_else_and_cse = PECoreRun_wen & mux_29_nl;
  assign and_1619_cse = while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1;
  assign nor_715_nl = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_2 | (~ or_dcpl_221));
  assign mux_545_nl = MUX_s_1_2_2(or_dcpl_221, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_546_nl = MUX_s_1_2_2(nor_715_nl, mux_545_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_547_nl = MUX_s_1_2_2(or_dcpl_221, mux_546_nl, while_stage_0_6);
  assign nor_716_nl = ~((~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1);
  assign mux_544_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_2, nor_716_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign nand_68_nl = ~(while_stage_0_6 & mux_544_nl);
  assign mux_548_nl = MUX_s_1_2_2(mux_547_nl, nand_68_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign mux_549_nl = MUX_s_1_2_2(and_1619_cse, mux_548_nl, nor_12_cse);
  assign and_1415_cse = mux_549_nl & PECoreRun_wen;
  assign weight_mem_banks_load_store_for_else_and_1_cse = PECoreRun_wen & and_1619_cse;
  assign weight_mem_banks_load_store_for_else_and_51_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign weight_mem_banks_load_store_for_else_and_53_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_mem_banks_load_store_for_else_and_54_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_mem_banks_load_store_for_else_and_57_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_mem_banks_load_store_for_else_and_59_cse = PECoreRun_wen & and_dcpl_48
      & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]))
      & nor_436_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign weight_mem_banks_load_store_for_else_and_62_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_247_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[23:16]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_247_nl);
  assign weight_read_addrs_and_17_cse = PECoreRun_wen & weight_mem_run_3_for_land_3_lpi_1_dfm_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign weight_read_addrs_and_19_cse = PECoreRun_wen & and_dcpl_90;
  assign weight_read_addrs_and_21_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse
      & and_dcpl_260;
  assign and_801_cse = (reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign and_802_cse = (reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2 | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign and_770_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1;
  assign and_776_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  assign and_771_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  assign and_773_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  assign and_774_cse = (reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign and_766_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  assign and_740_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1;
  assign and_767_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_3_sva;
  assign and_738_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  assign and_768_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  assign and_769_cse = (Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6 |
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign and_803_cse = (Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 |
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign and_804_cse = (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 |
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
      = weight_mem_read_arbxbar_arbiters_next_and_cse & or_dcpl_75;
  assign weight_read_addrs_and_30_enex5 = weight_write_data_data_and_16_cse & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  assign operator_15_false_1_and_cse = PECoreRun_wen & (~(and_113_cse | or_dcpl_75));
  assign PEManager_15U_PEManagerWrite_and_enex5 = PECoreRun_wen & reg_rva_in_reg_rw_sva_st_1_1_cse
      & (~ PECore_DecodeAxiWrite_switch_lp_nor_tmp_1) & PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1
      & (~ PECore_DecodeAxiWrite_switch_lp_equal_tmp_2) & (~ PECore_DecodeAxiWrite_switch_lp_equal_tmp_1)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_in_reg_data_sva_1_enexo;
  assign pe_manager_num_input_and_cse = PECoreRun_wen & (~(or_dcpl_249 | nand_88_cse
      | or_dcpl_284));
  assign pe_config_is_valid_and_cse = PECoreRun_wen & (~(PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1
      | PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (~ nand_88_cse);
  assign nor_721_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:10]!=2'b00));
  assign while_if_and_15_cse = PECoreRun_wen & and_dcpl_220;
  assign rva_in_reg_rw_and_6_cse = PECoreRun_wen & and_dcpl_83;
  assign rva_in_reg_rw_and_7_cse = PECoreRun_wen & and_dcpl_279;
  assign rva_in_reg_rw_and_8_cse = PECoreRun_wen & and_dcpl_280;
  assign while_if_and_16_cse = PECoreRun_wen & and_dcpl_281;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_398_cse = PECoreRun_wen
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp) & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_401_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_405_cse = PECoreRun_wen
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | weight_mem_run_3_for_weight_mem_run_3_for_and_1_tmp) & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_144_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_146_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_1_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign weight_port_read_out_data_and_174_cse = PECoreRun_wen & and_dcpl_280 & (~
      rva_in_reg_rw_sva_st_1_8) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  assign input_mem_banks_read_read_data_and_9_cse = PECoreRun_wen & and_dcpl_295
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6) & input_read_req_valid_lpi_1_dfm_1_8;
  assign weight_port_read_out_data_and_220_enex5 = weight_port_read_out_data_and_174_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo;
  assign input_mem_banks_read_read_data_and_51_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_52_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_53_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_54_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse = PECoreRun_wen & and_dcpl_280
      & (~(rva_in_reg_rw_sva_st_1_8 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6))
      & (~(input_read_req_valid_lpi_1_dfm_1_8 | rva_in_reg_rw_sva_8)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  assign PECore_RunMac_and_cse = (~ and_dcpl_24) & or_dcpl_287;
  assign PECore_RunMac_and_4_cse = and_dcpl_24 & or_dcpl_287;
  assign and_1446_cse = (PECore_UpdateFSM_switch_lp_equal_tmp_2_9 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
      | (~ while_stage_0_11) | (PECore_RunScale_PECore_RunScale_if_and_1_svs_8 &
      (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_8))) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & while_stage_0_10 & (PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8
      | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8));
  assign input_mem_banks_read_1_read_data_and_2_enex5 = PECoreRun_wen & PECore_RunMac_PECore_RunMac_if_and_svs_st_3
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  assign input_read_req_valid_and_1_cse = PECoreRun_wen & and_dcpl_295;
  assign PECore_DecodeAxiRead_switch_lp_and_7_cse = PECoreRun_wen & and_dcpl_308;
  assign rva_out_reg_data_and_40_cse = PECoreRun_wen & and_dcpl_308 & (~(rva_in_reg_rw_sva_st_8
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8))
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_8);
  assign rva_out_reg_data_and_157_enex5 = rva_out_reg_data_and_40_cse & reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_158_enex5 = rva_out_reg_data_and_40_cse & reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_159_enex5 = rva_out_reg_data_and_40_cse & reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  assign rva_out_reg_data_and_160_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_161_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_162_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_163_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_164_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_127_120_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_165_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_166_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_167_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_79_72_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_168_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_71_64_sva_dfm_4_3_enexo;
  assign ProductSum_for_and_cse = PECoreRun_wen & (or_dcpl_160 | and_dcpl_314);
  assign ProductSum_for_and_8_cse = (~ or_dcpl_160) & fsm_output;
  assign and_1462_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & while_stage_0_10;
  assign and_1464_cse = ((~((~(while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)))
      & fsm_output)) | and_1462_cse) & PECoreRun_wen;
  assign ProductSum_for_and_2_cse = PECoreRun_wen & and_1462_cse & and_dcpl_314;
  assign weight_port_read_out_data_and_182_ssc = PECoreRun_wen & and_dcpl_29 & (~
      rva_in_reg_rw_sva_st_1_7) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  assign weight_port_read_out_data_and_221_enex5 = weight_port_read_out_data_and_182_ssc
      & reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  assign weight_port_read_out_data_and_222_enex5 = weight_port_read_out_data_and_182_ssc
      & reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo;
  assign and_1476_cse = (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | PECore_UpdateFSM_switch_lp_equal_tmp_2_8)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & while_if_and_6_cse;
  assign PECore_RunScale_if_and_3_cse = PECoreRun_wen & and_dcpl_30;
  assign weight_mem_write_arbxbar_xbar_for_empty_and_enex5 = rva_in_reg_rw_and_6_cse
      & reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  assign and_319_cse = PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]);
  assign rva_in_reg_rw_and_11_cse = PECoreRun_wen & and_dcpl_41;
  assign pe_manager_base_weight_and_6_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse
      & and_dcpl_260;
  assign pe_manager_base_weight_and_7_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_3_or_cse
      & and_dcpl_260;
  assign input_mem_banks_read_read_data_and_18_cse = PECoreRun_wen & and_dcpl_346
      & input_read_req_valid_lpi_1_dfm_1_7 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5);
  assign input_mem_banks_read_read_data_and_55_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_56_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_57_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_58_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse = PECoreRun_wen & and_dcpl_351
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & (~ rva_in_reg_rw_sva_st_1_7) & (~(input_read_req_valid_lpi_1_dfm_1_7 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5))
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
  assign input_mem_banks_read_1_read_data_and_3_enex5 = PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_2 & while_stage_0_4 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  assign input_read_req_valid_and_2_cse = PECoreRun_wen & and_dcpl_346;
  assign PECore_DecodeAxiRead_switch_lp_and_11_cse = PECoreRun_wen & and_dcpl_359;
  assign rva_out_reg_data_and_58_cse = PECoreRun_wen & and_dcpl_359 & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_7 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7))
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 & (~ rva_in_reg_rw_sva_st_7);
  assign rva_out_reg_data_and_169_enex5 = rva_out_reg_data_and_58_cse & reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_170_enex5 = rva_out_reg_data_and_58_cse & reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_171_enex5 = rva_out_reg_data_and_58_cse & reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  assign weight_port_read_out_data_and_223_enex5 = weight_port_read_out_data_and_182_ssc
      & reg_weight_port_read_out_data_0_3_sva_dfm_2_enexo;
  assign weight_port_read_out_data_and_224_enex5 = weight_port_read_out_data_and_182_ssc
      & reg_weight_port_read_out_data_0_3_sva_dfm_2_1_enexo;
  assign rva_out_reg_data_and_172_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_173_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_174_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_175_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_176_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_127_120_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_177_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_119_112_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_178_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_111_104_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_179_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_180_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_79_72_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_181_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_71_64_sva_dfm_4_2_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_3_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp;
  assign PECore_RunMac_if_and_6_cse = PECoreRun_wen & and_666_cse;
  assign input_mem_banks_read_read_data_and_27_cse = PECoreRun_wen & and_dcpl_370
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4) & input_read_req_valid_lpi_1_dfm_1_6;
  assign input_mem_banks_read_read_data_and_59_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_60_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo;
  assign input_mem_banks_read_read_data_and_61_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_62_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse = PECoreRun_wen & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5
      & while_stage_0_8 & and_dcpl_374 & and_dcpl_373;
  assign and_380_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & PECore_UpdateFSM_switch_lp_equal_tmp_3_1 & while_stage_0_3;
  assign input_read_req_valid_and_3_cse = PECoreRun_wen & and_dcpl_370;
  assign PECore_DecodeAxiRead_switch_lp_and_15_cse = PECoreRun_wen & and_dcpl_370
      & and_dcpl_373;
  assign rva_out_reg_data_and_74_cse = PECoreRun_wen & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_6
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6))
      & (~ rva_in_reg_rw_sva_st_6) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5
      & while_stage_0_8 & and_dcpl_374 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4)
      & (~(rva_in_reg_rw_sva_6 | input_read_req_valid_lpi_1_dfm_1_6));
  assign rva_out_reg_data_and_182_enex5 = rva_out_reg_data_and_74_cse & reg_rva_out_reg_data_30_25_sva_dfm_4_enexo;
  assign rva_out_reg_data_and_183_enex5 = rva_out_reg_data_and_74_cse & reg_rva_out_reg_data_23_17_sva_dfm_4_enexo;
  assign rva_out_reg_data_and_184_enex5 = rva_out_reg_data_and_74_cse & reg_rva_out_reg_data_15_9_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_185_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_186_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_187_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_188_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_189_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_127_120_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_190_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_79_72_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_191_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_71_64_sva_dfm_4_1_enexo;
  assign PECore_RunScale_if_and_6_cse = PECoreRun_wen & and_dcpl_277;
  assign input_mem_banks_read_read_data_and_36_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      & while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~(rva_in_reg_rw_sva_st_1_5 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3));
  assign input_mem_banks_read_read_data_and_63_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  assign input_mem_banks_read_read_data_and_64_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1;
  assign input_mem_banks_read_read_data_and_65_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse = PECoreRun_wen & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1) & and_dcpl_41
      & and_dcpl_399;
  assign input_read_req_valid_and_4_cse = PECoreRun_wen & and_dcpl_403;
  assign PECore_DecodeAxiRead_switch_lp_and_19_cse = PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1)
      & while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & and_dcpl_399;
  assign rva_out_reg_data_and_90_cse = PECoreRun_wen & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_5)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5)
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      | rva_in_reg_rw_sva_st_5)) & and_dcpl_403 & (~(rva_in_reg_rw_sva_5 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3));
  assign rva_out_reg_data_and_192_enex5 = rva_out_reg_data_and_90_cse & reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_1_enexo;
  assign rva_out_reg_data_and_193_enex5 = rva_out_reg_data_and_90_cse & reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_1_enexo;
  assign rva_out_reg_data_and_194_enex5 = rva_out_reg_data_and_90_cse & reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_1_enexo;
  assign rva_out_reg_data_and_93_cse = PECoreRun_wen & and_dcpl_41 & (~(rva_in_reg_rw_sva_st_1_5
      & rva_in_reg_rw_sva_5));
  assign and_1489_cse = (~(((~(rva_in_reg_rw_sva_6 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      | (~ while_stage_0_8) | or_306_cse)) | rva_in_reg_rw_sva_st_1_5) & rva_in_reg_rw_sva_5))
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & PECoreRun_wen & while_stage_0_7;
  assign nor_462_nl = ~(rva_in_reg_rw_sva_st_1_5 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5));
  assign mux_96_nl = MUX_s_1_2_2(nor_462_nl, nand_32_cse, PECore_RunMac_PECore_RunMac_if_and_svs_st_5);
  assign rva_out_reg_data_and_98_cse = PECoreRun_wen & mux_96_nl & while_stage_0_7;
  assign PECore_RunScale_if_and_7_cse = PECoreRun_wen & and_dcpl_33;
  assign rva_out_reg_data_and_106_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (nand_40_cse | rva_in_reg_rw_sva_5);
  assign and_1506_cse = and_dcpl_279 & (~ rva_in_reg_rw_sva_6) & fsm_output & (rva_in_reg_rw_sva_5
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      | (~ while_stage_0_7)) & PECoreRun_wen;
  assign mux_33_nl = MUX_s_1_2_2((~ or_tmp_47), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign rva_out_reg_data_and_111_cse = PECoreRun_wen & mux_33_nl & and_dcpl_48;
  assign mux_101_nl = MUX_s_1_2_2(or_1109_cse, or_1106_cse, while_stage_0_5);
  assign mux_99_nl = MUX_s_1_2_2(reg_rva_in_reg_rw_sva_st_1_1_cse, or_1106_cse, while_stage_0_5);
  assign mux_100_nl = MUX_s_1_2_2(or_tmp_115, mux_99_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_102_nl = MUX_s_1_2_2(mux_101_nl, mux_100_nl, while_stage_0_3);
  assign mux_97_nl = MUX_s_1_2_2(reg_rva_in_reg_rw_sva_2_cse, or_1106_cse, while_stage_0_5);
  assign mux_98_nl = MUX_s_1_2_2(or_tmp_115, mux_97_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign mux_103_nl = MUX_s_1_2_2(mux_102_nl, mux_98_nl, while_stage_0_4);
  assign mux_104_nl = MUX_s_1_2_2(mux_103_nl, or_1105_cse, while_stage_0_6);
  assign rva_out_reg_data_and_112_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7 & fsm_output & mux_104_nl;
  assign nand_88_cse = ~(rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse);
  assign or_1106_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | rva_in_reg_rw_sva_3;
  assign or_1105_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | rva_in_reg_rw_sva_4;
  assign or_1109_cse = rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | nand_88_cse;
  assign or_1108_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign mux_551_nl = MUX_s_1_2_2(or_1109_cse, or_1108_nl, while_stage_0_3);
  assign or_1107_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | reg_rva_in_reg_rw_sva_2_cse;
  assign mux_552_nl = MUX_s_1_2_2(mux_551_nl, or_1107_nl, while_stage_0_4);
  assign mux_553_nl = MUX_s_1_2_2(mux_552_nl, or_1106_cse, while_stage_0_5);
  assign mux_554_nl = MUX_s_1_2_2(mux_553_nl, or_1105_cse, while_stage_0_6);
  assign and_1526_cse = mux_554_nl & fsm_output & while_stage_0_7 & PECoreRun_wen
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~ rva_in_reg_rw_sva_5);
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse = PECoreRun_wen & (~(rva_in_reg_rw_sva_st_1_4
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3
      & (~ rva_in_reg_rw_sva_4) & and_dcpl_48 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_106_nl = MUX_s_1_2_2((~ weight_mem_run_3_for_land_6_lpi_1_dfm_1), or_tmp_47,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_107_nl = MUX_s_1_2_2(mux_106_nl, or_tmp_7, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign PECore_DecodeAxiRead_switch_lp_and_23_cse = PECoreRun_wen & (~ mux_107_nl)
      & while_stage_0_6;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_24_cse = PECoreRun_wen & and_dcpl_435
      & and_dcpl_434 & and_dcpl_433;
  assign input_mem_banks_read_read_data_and_45_enex5 = PECoreRun_wen & and_dcpl_435
      & input_read_req_valid_lpi_1_dfm_1_3 & and_dcpl_83 & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo;
  assign nor_465_nl = ~(rva_in_reg_rw_sva_3 | input_read_req_valid_lpi_1_dfm_1_3
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1);
  assign mux_109_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, nor_465_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign PECore_DecodeAxiRead_switch_lp_and_27_cse = PECoreRun_wen & mux_109_nl &
      while_stage_0_5;
  assign rva_out_reg_data_and_120_cse = PECoreRun_wen & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_3
      | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1))
      & and_dcpl_434 & (~ rva_in_reg_rw_sva_3) & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 | rva_in_reg_rw_sva_st_3)) &
      and_dcpl_83;
  assign rva_out_reg_data_and_195_enex5 = rva_out_reg_data_and_120_cse & reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_196_enex5 = rva_out_reg_data_and_120_cse & reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_197_enex5 = rva_out_reg_data_and_120_cse & reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_123_cse = PECoreRun_wen & and_dcpl_435 & (~ input_read_req_valid_lpi_1_dfm_1_3)
      & and_dcpl_433;
  assign rva_out_reg_data_and_198_enex5 = rva_out_reg_data_and_123_cse & reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_199_enex5 = rva_out_reg_data_and_123_cse & reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_200_enex5 = rva_out_reg_data_and_123_cse & reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_201_enex5 = rva_out_reg_data_and_123_cse & reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_202_enex5 = rva_out_reg_data_and_123_cse & reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_29_cse = PECoreRun_wen & and_dcpl_458
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 & and_dcpl_172;
  assign input_mem_banks_read_read_data_and_46_enex5 = PECoreRun_wen & or_dcpl_201
      & (~ reg_rva_in_reg_rw_sva_2_cse) & input_read_req_valid_lpi_1_dfm_1_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1;
  assign PECore_DecodeAxiRead_switch_lp_and_31_cse = PECoreRun_wen & and_dcpl_458
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign rva_out_reg_data_and_128_cse = PECoreRun_wen & (~(input_read_req_valid_lpi_1_dfm_1_2
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_2)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2))
      & (~ reg_rva_in_reg_rw_sva_2_cse) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign rva_out_reg_data_and_203_enex5 = rva_out_reg_data_and_128_cse & reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  assign rva_out_reg_data_and_204_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_205_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_206_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_207_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_208_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse = PECoreRun_wen & mux_tmp_110
      & and_dcpl_480;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_35_cse = PECoreRun_wen & (~ reg_rva_in_reg_rw_sva_st_1_1_cse)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_switch_lp_and_35_cse = PECoreRun_wen & and_dcpl_480;
  assign rva_out_reg_data_and_136_enex5 = PECoreRun_wen & (~(input_read_req_valid_lpi_1_dfm_1_1
      | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[0])))
      & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[3:1]==3'b010)
      & and_dcpl_488 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_209_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_210_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_211_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_212_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_213_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_pe_config_input_counter_sva_dfm_1_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse = PECoreRun_wen & mux_tmp_110
      & and_dcpl_479 & (~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1) &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse = PECoreRun_wen & and_dcpl_227
      & reg_rva_in_PopNB_mioi_iswt0_cse & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))
      & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_44_cse = PECoreRun_wen & and_dcpl_321
      & and_dcpl_220 & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt))
      & nand_41_cse;
  assign rva_out_reg_data_and_143_cse = PECoreRun_wen & ((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]!=4'b0110))
      & and_dcpl_281;
  assign and_568_cse = while_stage_0_12 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
      & (~ rva_in_reg_rw_sva_st_1_10);
  assign or_380_cse = (state_2_1_sva!=2'b00) | state_0_sva;
  assign weight_mem_run_3_for_5_and_145_cse = reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_port_read_out_data_0_7_sva_mx0 = MUX1HOT_v_8_3_2(({weight_port_read_out_data_0_3_sva_dfm_1_1_7_4
      , weight_port_read_out_data_0_3_sva_dfm_1_1_3_0}), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1,
      weight_port_read_out_data_0_7_sva, {and_dcpl_279 , and_dcpl_277 , (~ while_stage_0_8)});
  assign PECore_PushAxiRsp_if_else_mux_23_mx0w2 = MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1);
  assign mux1h_4_nl = MUX1HOT_v_8_7_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[63:56]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63:56]),
      weight_port_read_out_data_0_7_sva_mx0, {and_1147_cse , and_1148_cse , and_1149_cse
      , and_1150_cse , and_1151_cse , and_1152_cse , nor_626_cse});
  assign not_2376_nl = ~ or_dcpl;
  assign weight_port_read_out_data_0_7_sva_dfm_mx0w2 = MUX_v_8_2_2(8'b00000000, mux1h_4_nl,
      not_2376_nl);
  assign or_894_tmp = ((pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2) | and_dcpl;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign Arbiter_8U_Roundrobin_pick_nand_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1)
      & and_dcpl_90)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_38_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1
      & and_dcpl_90;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_56_nl = weight_mem_read_arbxbar_arbiters_next_7_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_56_nl,
      weight_mem_read_arbxbar_arbiters_next_7_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_57_nl = weight_mem_read_arbxbar_arbiters_next_7_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_57_nl,
      weight_mem_read_arbxbar_arbiters_next_7_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_58_nl = weight_mem_read_arbxbar_arbiters_next_7_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_58_nl,
      weight_mem_read_arbxbar_arbiters_next_7_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_59_nl = weight_mem_read_arbxbar_arbiters_next_7_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_59_nl,
      weight_mem_read_arbxbar_arbiters_next_7_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_60_nl = weight_mem_read_arbxbar_arbiters_next_7_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_60_nl,
      weight_mem_read_arbxbar_arbiters_next_7_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_61_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_61_nl,
      weight_mem_read_arbxbar_arbiters_next_7_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_90);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign Arbiter_8U_Roundrobin_pick_nand_42_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)
      & and_dcpl_90)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_37_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1
      & and_dcpl_90;
  assign weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_90);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign Arbiter_8U_Roundrobin_pick_1_mux_429_mx1w1 = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign Arbiter_8U_Roundrobin_pick_or_3_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1)
      & and_dcpl_90)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_7_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1
      & and_dcpl_90;
  assign weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_3_cse , Arbiter_8U_Roundrobin_pick_and_7_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign Arbiter_8U_Roundrobin_pick_1_mux_428_mx1w1 = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_3_cse , Arbiter_8U_Roundrobin_pick_and_7_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl = weight_mem_read_arbxbar_arbiters_next_5_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl,
      weight_mem_read_arbxbar_arbiters_next_5_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_3_cse , Arbiter_8U_Roundrobin_pick_and_7_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl = weight_mem_read_arbxbar_arbiters_next_5_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl,
      weight_mem_read_arbxbar_arbiters_next_5_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_3_cse , Arbiter_8U_Roundrobin_pick_and_7_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_nl = weight_mem_read_arbxbar_arbiters_next_5_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_nl,
      weight_mem_read_arbxbar_arbiters_next_5_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_3_cse , Arbiter_8U_Roundrobin_pick_and_7_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_73_nl = weight_mem_read_arbxbar_arbiters_next_5_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_73_nl,
      weight_mem_read_arbxbar_arbiters_next_5_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_3_cse , Arbiter_8U_Roundrobin_pick_and_7_cse});
  assign weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_90);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign Arbiter_8U_Roundrobin_pick_nand_30_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1)
      & and_dcpl_90)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_31_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1
      & and_dcpl_90;
  assign weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_33_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_33_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_90);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign Arbiter_8U_Roundrobin_pick_nand_18_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1)
      & and_dcpl_90)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_25_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1
      & and_dcpl_90;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_83_nl = weight_mem_read_arbxbar_arbiters_next_3_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_83_nl,
      weight_mem_read_arbxbar_arbiters_next_3_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_90);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_20_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign Arbiter_8U_Roundrobin_pick_nand_8_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1)
      & and_dcpl_90)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_20_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1
      & and_dcpl_90;
  assign weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_20_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_19_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_19_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_18_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_18_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_17_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_17_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl,
      weight_mem_read_arbxbar_arbiters_next_2_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_15_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_15_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_90);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign Arbiter_8U_Roundrobin_pick_or_1_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1)
      & and_dcpl_90)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_3_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1
      & and_dcpl_90;
  assign weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_1_cse , Arbiter_8U_Roundrobin_pick_and_3_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl = weight_mem_read_arbxbar_arbiters_next_1_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl,
      weight_mem_read_arbxbar_arbiters_next_1_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_1_cse , Arbiter_8U_Roundrobin_pick_and_3_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl = weight_mem_read_arbxbar_arbiters_next_1_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl,
      weight_mem_read_arbxbar_arbiters_next_1_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_1_cse , Arbiter_8U_Roundrobin_pick_and_3_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_1_cse , Arbiter_8U_Roundrobin_pick_and_3_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl,
      weight_mem_read_arbxbar_arbiters_next_1_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_1_cse , Arbiter_8U_Roundrobin_pick_and_3_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_nl,
      weight_mem_read_arbxbar_arbiters_next_1_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_or_1_cse , Arbiter_8U_Roundrobin_pick_and_3_cse});
  assign weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_90);
  assign Arbiter_8U_Roundrobin_pick_nand_77_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1)
      & and_dcpl_90)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_54_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1
      & and_dcpl_90;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_98_nl = weight_mem_read_arbxbar_arbiters_next_0_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_98_nl,
      weight_mem_read_arbxbar_arbiters_next_0_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_77_cse , Arbiter_8U_Roundrobin_pick_and_54_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_99_nl = weight_mem_read_arbxbar_arbiters_next_0_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_99_nl,
      weight_mem_read_arbxbar_arbiters_next_0_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_77_cse , Arbiter_8U_Roundrobin_pick_and_54_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl = weight_mem_read_arbxbar_arbiters_next_0_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl,
      weight_mem_read_arbxbar_arbiters_next_0_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_77_cse , Arbiter_8U_Roundrobin_pick_and_54_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl = weight_mem_read_arbxbar_arbiters_next_0_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl,
      weight_mem_read_arbxbar_arbiters_next_0_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_77_cse , Arbiter_8U_Roundrobin_pick_and_54_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl = weight_mem_read_arbxbar_arbiters_next_0_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl,
      weight_mem_read_arbxbar_arbiters_next_0_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_77_cse , Arbiter_8U_Roundrobin_pick_and_54_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_103_nl = weight_mem_read_arbxbar_arbiters_next_0_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_103_nl,
      weight_mem_read_arbxbar_arbiters_next_0_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1,
      {and_dcpl_83 , Arbiter_8U_Roundrobin_pick_nand_77_cse , Arbiter_8U_Roundrobin_pick_and_54_cse});
  assign weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_90);
  assign pe_manager_base_weight_sva_mx1_3_0 = MUX_v_4_2_2((pe_manager_base_weight_sva[3:0]),
      (pe_manager_base_weight_sva_dfm_3_1[3:0]), while_stage_0_5);
  assign pe_manager_base_weight_sva_mx2 = MUX_v_15_2_2(pe_manager_base_weight_sva,
      pe_manager_base_weight_sva_dfm_3_1, while_stage_0_5);
  assign pe_manager_base_weight_sva_mx3_0 = MUX_s_1_2_2((pe_manager_base_weight_sva[0]),
      (pe_manager_base_weight_sva_dfm_3_1[0]), while_stage_0_5);
  assign nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000001;
  assign PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_1_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000001;
  assign operator_15_false_acc_nl = nl_operator_15_false_acc_nl[13:0];
  assign weight_read_addrs_2_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000011;
  assign PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_3_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_1_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:2])}) + 13'b0000000000001;
  assign operator_15_false_acc_1_nl = nl_operator_15_false_acc_1_nl[12:0];
  assign weight_read_addrs_4_14_2_lpi_1_dfm_1_1 = MUX_v_13_2_2(13'b0000000000000,
      operator_15_false_acc_1_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000101;
  assign PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_5_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_2_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000011;
  assign operator_15_false_acc_2_nl = nl_operator_15_false_acc_2_nl[13:0];
  assign weight_read_addrs_6_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_2_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000111;
  assign PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_7_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112, and_113_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97, and_120_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82, and_127_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67, and_134_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52, and_141_cse);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_15_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37, and_148_cse);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22, and_dcpl_643);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7, and_162_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1 = (state_2_1_sva[0]) & (~((state_2_1_sva[1])
      | state_0_sva));
  assign state_mux_1_cse = MUX_v_2_2_2(state_2_1_sva, state_2_1_sva_dfm_1, while_stage_0_3);
  assign state_0_sva_mx1 = MUX_s_1_2_2(PECore_UpdateFSM_next_state_0_lpi_1_dfm_4,
      state_0_sva, or_dcpl_237);
  assign pe_config_manager_counter_sva_mx1 = MUX_v_4_2_2(pe_config_manager_counter_sva,
      pe_config_manager_counter_sva_dfm_3_1, and_1341_cse);
  assign PECore_PushOutput_PECore_PushOutput_if_and_svs_1 = (state_mux_1_cse[1])
      & (~((state_mux_1_cse[0]) | state_0_sva_mx1));
  assign PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1 = ~(PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_380_cse);
  assign pe_config_input_counter_and_cse = while_if_and_tmp_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign nl_operator_8_false_acc_nl = pe_config_input_counter_sva + 8'b00000001;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[7:0];
  assign pe_config_UpdateInputCounter_not_nl = ~ pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl = MUX_v_8_2_2(8'b00000000,
      operator_8_false_acc_nl, pe_config_UpdateInputCounter_not_nl);
  assign pe_config_input_counter_nand_nl = ~(while_stage_0_3 & (~((~(PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1266_cse_1)));
  assign pe_config_input_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_input_counter_sva,
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl, pe_config_input_counter_sva_dfm_1,
      {pe_config_input_counter_nand_nl , and_380_cse , pe_config_input_counter_and_cse});
  assign nl_operator_8_false_1_acc_nl = pe_config_output_counter_sva + 8'b00000001;
  assign operator_8_false_1_acc_nl = nl_operator_8_false_1_acc_nl[7:0];
  assign pe_config_UpdateManagerCounter_if_not_9_nl = ~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl
      = MUX_v_8_2_2(8'b00000000, operator_8_false_1_acc_nl, pe_config_UpdateManagerCounter_if_not_9_nl);
  assign pe_config_output_counter_nand_nl = ~(while_stage_0_3 & (~((~(PECore_UpdateFSM_switch_lp_and_2_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1266_cse_1)));
  assign while_and_152_nl = PECore_UpdateFSM_switch_lp_and_2_tmp_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign pe_config_output_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_output_counter_sva,
      pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl,
      pe_config_output_counter_sva_dfm_1, {pe_config_output_counter_nand_nl , while_and_152_nl
      , pe_config_input_counter_and_cse});
  assign and_666_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_if_and_2_m1c = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & and_666_cse;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl
      = pe_config_is_zero_first_sva & (~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1);
  assign while_if_or_nl = (~((~((~ PECore_UpdateFSM_switch_lp_equal_tmp_5_1) & and_666_cse))
      & while_stage_0_3)) | ((~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1)
      & while_if_and_2_m1c);
  assign while_if_and_4_nl = pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
      & while_if_and_2_m1c;
  assign pe_config_is_zero_first_sva_mx1 = MUX1HOT_s_1_3_2(while_if_mux_27_itm_1,
      pe_config_is_zero_first_sva, pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl,
      {and_dcpl_212 , while_if_or_nl , while_if_and_4_nl});
  assign PECore_UpdateFSM_switch_lp_equal_tmp_6 = state_0_sva_mx1 & (state_mux_1_cse==2'b00);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1 = (state_mux_1_cse[0])
      & (~((state_mux_1_cse[1]) | state_0_sva_mx1));
  assign pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1
      = ~((pe_config_manager_counter_sva_mx1 != (operator_4_false_acc_sdt_sva_1[3:0]))
      | (operator_4_false_acc_sdt_sva_1[4]));
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0110);
  assign PECore_UpdateFSM_switch_lp_not_27_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_nl
      = MUX_v_17_2_2(17'b00000000000000000, act_port_reg_data_48_32_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_27_nl);
  assign act_port_reg_data_48_32_sva_mx1 = MUX_v_17_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_nl,
      act_port_reg_data_48_32_sva, or_dcpl_257);
  assign PECore_UpdateFSM_switch_lp_not_28_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_nl
      = MUX_v_17_2_2(17'b00000000000000000, act_port_reg_data_80_64_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_28_nl);
  assign act_port_reg_data_80_64_sva_mx1 = MUX_v_17_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_nl,
      act_port_reg_data_80_64_sva, or_dcpl_257);
  assign PECore_UpdateFSM_switch_lp_not_29_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_nl
      = MUX_v_17_2_2(17'b00000000000000000, act_port_reg_data_112_96_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_29_nl);
  assign act_port_reg_data_112_96_sva_mx1 = MUX_v_17_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_nl,
      act_port_reg_data_112_96_sva, or_dcpl_257);
  assign PECore_UpdateFSM_switch_lp_not_19_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_11_nl
      = MUX_v_17_2_2(17'b00000000000000000, act_port_reg_data_144_128_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_19_nl);
  assign act_port_reg_data_144_128_sva_mx1 = MUX_v_17_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_11_nl,
      act_port_reg_data_144_128_sva, or_dcpl_257);
  assign weight_mem_run_3_for_weight_mem_run_3_for_and_7_tmp = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1);
  assign weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1);
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp;
  assign weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse;
  assign weight_mem_run_3_for_weight_mem_run_3_for_and_1_tmp = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6,
      or_dcpl_236);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0,
      or_dcpl_236);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5,
      or_dcpl_236);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1,
      or_dcpl_236);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4,
      or_dcpl_236);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2,
      or_dcpl_236);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3,
      or_dcpl_236);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0101);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b111)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1 = (pe_manager_base_weight_sva[2:0]==3'b110)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b100)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b010)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b001)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign weight_mem_run_3_for_weight_mem_run_3_for_and_6_tmp = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_1);
  assign weight_mem_run_3_for_land_1_lpi_1_dfm_1_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_15_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1 = MUX_v_3_2_2(3'b000,
      (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0]), weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp = MUX_s_1_8_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp
      | (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp));
  assign while_and_221_rgt = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_225_rgt = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_229_rgt = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_233_rgt = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_237_rgt = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_241_rgt = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_245_rgt = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_249_rgt = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_253_rgt = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_257_rgt = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_261_rgt = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_265_rgt = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_269_rgt = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_273_rgt = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_277_rgt = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_281_rgt = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_285_rgt = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_289_rgt = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_293_rgt = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_297_rgt = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_301_rgt = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_305_rgt = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_309_rgt = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_313_rgt = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_317_rgt = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_321_rgt = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_325_rgt = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_329_rgt = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_333_rgt = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_337_rgt = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_341_rgt = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_345_rgt = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_349_rgt = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_353_rgt = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_357_rgt = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_361_rgt = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_365_rgt = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_369_rgt = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_373_rgt = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_377_rgt = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_381_rgt = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_385_rgt = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_389_rgt = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_393_rgt = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_397_rgt = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_401_rgt = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_405_rgt = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_409_rgt = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_413_rgt = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_417_rgt = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_421_rgt = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_425_rgt = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_429_rgt = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_433_rgt = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_437_rgt = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_441_rgt = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_445_rgt = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_449_rgt = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_453_rgt = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_457_rgt = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_461_rgt = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_465_rgt = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_469_rgt = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_473_rgt = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_477_rgt = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_481_rgt = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_485_rgt = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_489_rgt = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_493_rgt = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_497_rgt = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_501_rgt = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_505_rgt = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_509_rgt = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_513_rgt = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_517_rgt = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_521_rgt = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_525_rgt = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_529_rgt = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_533_rgt = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_537_rgt = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_541_rgt = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_545_rgt = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_549_rgt = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_553_rgt = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_557_rgt = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_561_rgt = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_565_rgt = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_569_rgt = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_573_rgt = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_577_rgt = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_581_rgt = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_585_rgt = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_589_rgt = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_593_rgt = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_597_rgt = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_601_rgt = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_605_rgt = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_609_rgt = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_613_rgt = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_617_rgt = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_621_rgt = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_625_rgt = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_629_rgt = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_633_rgt = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_637_rgt = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_641_rgt = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_645_rgt = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_649_rgt = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_653_rgt = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_657_rgt = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_661_rgt = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_665_rgt = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_669_rgt = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_673_rgt = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_677_rgt = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_681_rgt = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_685_rgt = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_689_rgt = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_693_rgt = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_697_rgt = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_701_rgt = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_705_rgt = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_709_rgt = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_713_rgt = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_717_rgt = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_721_rgt = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_725_rgt = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_729_rgt = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_733_rgt = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_737_rgt = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_741_rgt = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_745_rgt = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_749_rgt = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_753_rgt = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_757_rgt = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_761_rgt = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_765_rgt = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_769_rgt = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_773_rgt = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_777_rgt = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_781_rgt = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_785_rgt = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_789_rgt = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_793_rgt = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_797_rgt = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_801_rgt = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_805_rgt = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_809_rgt = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_813_rgt = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_817_rgt = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_821_rgt = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_825_rgt = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_829_rgt = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_833_rgt = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_837_rgt = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_841_rgt = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_845_rgt = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_849_rgt = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_853_rgt = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_857_rgt = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_861_rgt = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_865_rgt = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_869_rgt = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_873_rgt = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_877_rgt = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_881_rgt = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_885_rgt = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_889_rgt = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_893_rgt = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_897_rgt = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_901_rgt = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_905_rgt = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_909_rgt = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_913_rgt = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_917_rgt = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_921_rgt = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_925_rgt = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_929_rgt = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_933_rgt = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_937_rgt = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_941_rgt = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_945_rgt = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_949_rgt = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_953_rgt = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_957_rgt = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_961_rgt = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_965_rgt = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_969_rgt = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_973_rgt = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_977_rgt = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_981_rgt = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_985_rgt = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_989_rgt = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_993_rgt = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_997_rgt = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1001_rgt = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1005_rgt = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1009_rgt = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1013_rgt = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1017_rgt = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1021_rgt = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1025_rgt = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1029_rgt = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1033_rgt = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1037_rgt = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1041_rgt = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1045_rgt = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1049_rgt = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1053_rgt = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1057_rgt = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1061_rgt = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1065_rgt = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1069_rgt = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1073_rgt = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1077_rgt = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1081_rgt = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1085_rgt = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1089_rgt = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1093_rgt = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1097_rgt = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1101_rgt = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1105_rgt = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1109_rgt = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1113_rgt = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1117_rgt = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1121_rgt = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1125_rgt = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1129_rgt = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1133_rgt = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1137_rgt = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1141_rgt = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1145_rgt = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1149_rgt = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1153_rgt = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1157_rgt = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1161_rgt = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1165_rgt = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1169_rgt = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1173_rgt = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1177_rgt = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1181_rgt = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1185_rgt = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1189_rgt = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1193_rgt = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1197_rgt = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1201_rgt = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1205_rgt = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1209_rgt = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1213_rgt = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1217_rgt = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1221_rgt = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1225_rgt = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1229_rgt = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1233_rgt = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1237_rgt = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1241_rgt = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign PECore_PushAxiRsp_mux_24_nl = MUX_s_1_2_2(reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse,
      PECore_PushAxiRsp_mux_10_itm_1, rva_in_reg_rw_sva_5);
  assign PECore_PushAxiRsp_if_else_mux_10_mx0w2 = MUX_s_1_2_2(PECore_PushAxiRsp_mux_24_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1);
  assign while_if_while_if_and_24_nl = MUX_v_8_2_2(8'b00000000, rva_out_reg_data_127_120_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_127_120_sva_dfm_4_mx0w0 = MUX1HOT_v_8_3_2(while_if_while_if_and_24_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_30_nl = MUX_v_8_2_2(8'b00000000, rva_out_reg_data_79_72_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_79_72_sva_dfm_7 = MUX1HOT_v_8_3_2(while_if_while_if_and_30_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_31_nl = MUX_v_8_2_2(8'b00000000, rva_out_reg_data_71_64_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_71_64_sva_dfm_7 = MUX1HOT_v_8_3_2(while_if_while_if_and_31_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_55_48_sva_dfm_6_mx1 = MUX_v_8_2_2(rva_out_reg_data_55_48_sva_dfm_4_1,
      rva_out_reg_data_55_48_sva_dfm_6, or_dcpl_291);
  assign rva_out_reg_data_62_56_sva_dfm_6_mx1 = MUX_v_7_2_2(rva_out_reg_data_62_56_sva_dfm_4_1,
      rva_out_reg_data_62_56_sva_dfm_6, or_dcpl_291);
  assign rva_out_reg_data_46_40_sva_dfm_6_mx1 = MUX_v_7_2_2(rva_out_reg_data_46_40_sva_dfm_4_1,
      rva_out_reg_data_46_40_sva_dfm_6, or_dcpl_291);
  assign rva_out_reg_data_35_32_sva_dfm_6_mx1 = MUX_v_4_2_2(rva_out_reg_data_35_32_sva_dfm_4_1,
      rva_out_reg_data_35_32_sva_dfm_6, or_dcpl_291);
  assign pe_manager_base_input_sva_mx1_7_0 = MUX_v_8_2_2((pe_manager_base_input_sva[7:0]),
      (pe_manager_base_input_sva_dfm_3_1[7:0]), while_stage_0_3);
  assign pe_manager_base_input_sva_mx2 = MUX_v_15_2_2(pe_manager_base_input_sva,
      pe_manager_base_input_sva_dfm_3_1, while_stage_0_3);
  assign PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
      & PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3
      | and_319_cse);
  assign PECore_RunScale_PECore_RunScale_if_and_1_svs_1 = (state_mux_1_cse[0]) &
      state_0_sva_mx1 & (~ (state_mux_1_cse[1]));
  assign PECore_DecodeAxiRead_switch_lp_nor_tmp_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_DecodeAxiRead_switch_lp_nor_9_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 | PECore_DecodeAxiRead_switch_lp_nor_tmp_10);
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1 = ~(input_read_req_valid_lpi_1_dfm_1_10
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse});
  assign weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0 = MUX_v_128_2_2(weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0 = MUX_v_120_2_2(weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_8,
      (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:8]), weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_load_store_1_for_else_else_and_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_or_nl = (weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1);
  assign weight_mem_banks_load_store_1_for_else_else_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9 = MUX1HOT_v_8_6_2(BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8,
      ({weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7
      , weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_6_0}),
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1,
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[7:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[7:0]),
      {weight_mem_banks_load_store_1_for_else_else_and_nl , weight_mem_banks_load_store_1_for_else_else_or_nl
      , weight_mem_banks_load_store_1_for_else_else_and_4_nl , weight_mem_banks_load_store_1_for_else_else_and_6_nl
      , weight_mem_banks_load_store_1_for_else_else_and_8_nl , weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {weight_mem_run_3_for_5_and_145_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_weight_mem_run_3_for_5_and_151_itm_2_cse , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {weight_mem_run_3_for_5_and_145_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_weight_mem_run_3_for_5_and_151_itm_2_cse , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {weight_mem_run_3_for_5_and_145_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_weight_mem_run_3_for_5_and_151_itm_2_cse , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {weight_mem_run_3_for_5_and_145_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_weight_mem_run_3_for_5_and_151_itm_2_cse , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {weight_mem_run_3_for_5_and_145_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_weight_mem_run_3_for_5_and_151_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {weight_mem_run_3_for_5_and_145_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_21_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_21_nl
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2_cse , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 , reg_weight_mem_run_3_for_5_and_151_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {weight_mem_run_3_for_5_and_145_cse
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 , reg_weight_mem_run_3_for_5_and_151_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_nl
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse = reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_14_itm_1_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_14_itm_1_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1
      , weight_mem_run_3_for_5_asn_459 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_265_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_265_nl , weight_mem_run_3_for_5_asn_455
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_4_itm_2_cse
      , weight_mem_run_3_for_5_asn_459 , reg_weight_mem_run_3_for_5_and_6_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1 , PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367
      , weight_mem_run_3_for_5_asn_455 , weight_mem_run_3_for_5_asn_457 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_2
      , weight_mem_run_3_for_5_asn_459 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_69_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_69_nl , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_weight_mem_run_3_for_5_and_151_itm_2_cse , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
      {weight_mem_run_3_for_5_and_145_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_2
      , reg_weight_mem_run_3_for_5_and_151_itm_2_cse , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
      {weight_mem_run_3_for_5_and_145_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_weight_mem_run_3_for_5_and_151_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
      {weight_mem_run_3_for_5_and_145_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
      {weight_mem_run_3_for_5_and_145_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
      {weight_mem_run_3_for_5_and_145_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , reg_weight_mem_run_3_for_5_and_151_itm_2_cse , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b100)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1 = (~(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_sva_1) & not_tmp_404;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_sva_1 & not_tmp_404;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_sva_1 | mux_192_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_sva_1 & (~ mux_192_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_sva_1) & and_dcpl_698;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_sva_1 & and_dcpl_698;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]),
      {mux_tmp_166 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_sva_1,
      {mux_tmp_166 , not_tmp_404 , (~ mux_192_itm) , and_dcpl_698});
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  assign mux_202_nl = MUX_s_1_2_2(mux_tmp_185, mux_tmp_183, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl,
      mux_202_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 | mux_214_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 & (~ mux_214_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 | mux_228_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 & (~ mux_228_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1) & and_dcpl_701;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 & and_dcpl_701;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]),
      {mux_tmp_205 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1,
      {mux_tmp_205 , (~ mux_214_itm) , (~ mux_228_itm) , and_dcpl_701});
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  assign mux_237_nl = MUX_s_1_2_2(or_tmp_270, or_tmp_265, while_stage_0_5);
  assign or_566_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | or_tmp_270;
  assign or_561_nl = while_mux_1438_tmp | or_tmp_265;
  assign mux_236_nl = MUX_s_1_2_2(or_566_nl, or_561_nl, while_stage_0_5);
  assign mux_238_nl = MUX_s_1_2_2(mux_237_nl, mux_236_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl,
      mux_238_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1) & not_tmp_417;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 & not_tmp_417;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1) & not_tmp_419;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 & not_tmp_419;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1) & and_dcpl_703;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 & and_dcpl_703;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]),
      {mux_tmp_244 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1,
      {mux_tmp_244 , not_tmp_417 , not_tmp_419 , and_dcpl_703});
  assign and_1100_cse = Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign and_1101_cse = Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign and_1092_cse = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign and_1094_cse = weight_mem_read_arbxbar_arbiters_next_5_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign and_1093_cse = weight_mem_read_arbxbar_arbiters_next_5_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign and_1095_cse = while_mux_1430_tmp & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign and_1098_cse = Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign while_mux_1435_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_428_mx1w1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_1097_cse = while_mux_1435_nl & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign while_mux_1436_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_429_mx1w1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_1096_cse = while_mux_1436_nl & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign and_1099_cse = Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign or_628_nl = and_1098_cse | and_1099_cse | and_1100_cse | and_1101_cse;
  assign mux_284_nl = MUX_s_1_2_2(or_tmp_287, or_628_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_622_nl = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign mux_283_nl = MUX_s_1_2_2(or_tmp_287, or_622_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign mux_285_cse = MUX_s_1_2_2(mux_284_nl, mux_283_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign nor_617_nl = ~(and_1092_cse | and_1093_cse | and_1094_cse | or_tmp_287);
  assign nor_618_nl = ~(and_1095_cse | and_1096_cse | and_1097_cse | mux_285_cse);
  assign mux_286_nl = MUX_s_1_2_2(nor_617_nl, nor_618_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl,
      mux_286_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 | mux_304_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 & (~ mux_304_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 | mux_322_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 & (~ mux_322_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1) & and_dcpl_706;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 & and_dcpl_706;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]),
      {mux_tmp_288 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1,
      {mux_tmp_288 , (~ mux_304_itm) , (~ mux_322_itm) , and_dcpl_706});
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1;
  assign mux_335_nl = MUX_s_1_2_2(or_tmp_395, or_tmp_389, while_stage_0_5);
  assign or_695_nl = weight_mem_read_arbxbar_arbiters_next_4_3_sva | or_tmp_395;
  assign or_694_nl = while_mux_1427_tmp | or_tmp_389;
  assign mux_334_nl = MUX_s_1_2_2(or_695_nl, or_694_nl, while_stage_0_5);
  assign mux_336_nl = MUX_s_1_2_2(mux_335_nl, mux_334_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign or_693_nl = weight_mem_read_arbxbar_arbiters_next_4_1_sva | or_tmp_395;
  assign or_692_nl = while_mux_1429_tmp | or_tmp_389;
  assign mux_332_nl = MUX_s_1_2_2(or_693_nl, or_692_nl, while_stage_0_5);
  assign or_691_nl = or_tmp_348 | or_tmp_395;
  assign or_685_nl = or_tmp_345 | or_tmp_389;
  assign mux_331_nl = MUX_s_1_2_2(or_691_nl, or_685_nl, while_stage_0_5);
  assign mux_333_nl = MUX_s_1_2_2(mux_332_nl, mux_331_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign mux_337_nl = MUX_s_1_2_2(mux_336_nl, mux_333_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl,
      mux_337_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_nl
      = weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 | mux_347_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 & (~ mux_347_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1) & and_dcpl_707;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 & and_dcpl_707;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1) & and_dcpl_712;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 & and_dcpl_712;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]),
      {mux_tmp_338 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1,
      {mux_tmp_338 , (~ mux_347_itm) , and_dcpl_707 , and_dcpl_712});
  assign and_1107_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) & while_mux_1417_tmp;
  assign and_1110_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]) & while_mux_1416_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_mux_608_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1421_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_608_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_1108_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) & while_mux_1421_nl;
  assign and_1106_cse = weight_mem_read_arbxbar_arbiters_next_3_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign and_1109_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]) & while_mux_1420_tmp;
  assign and_1111_cse = while_mux_1422_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign or_885_nl = and_771_cse | and_776_cse | and_773_cse | and_770_cse | and_1106_cse
      | and_789_cse;
  assign or_886_nl = and_1107_cse | and_1108_cse | and_1109_cse | and_1110_cse |
      and_1111_cse | nor_tmp_230;
  assign mux_362_nl = MUX_s_1_2_2(or_885_nl, or_886_nl, while_stage_0_5);
  assign nor_621_nl = ~(mux_362_nl | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl,
      nor_621_nl);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | (weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]));
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 | mux_387_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 & (~ mux_387_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_32_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1) & not_tmp_443;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 & not_tmp_443;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1) & and_dcpl_717;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 & and_dcpl_717;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]),
      {mux_tmp_366 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_32_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1,
      {mux_tmp_366 , (~ mux_387_itm) , not_tmp_443 , and_dcpl_717});
  assign and_1114_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  assign and_1118_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]) & while_mux_1413_tmp;
  assign and_1119_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) & while_mux_1414_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign nor_622_nl = ~(and_767_cse | and_738_cse | and_1114_cse | and_766_cse |
      and_740_cse | and_768_cse | and_1028_cse);
  assign or_794_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva | or_tmp_496;
  assign or_793_nl = Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 | or_tmp_496;
  assign mux_404_nl = MUX_s_1_2_2(or_794_nl, or_793_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_792_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2])
      | weight_mem_read_arbxbar_arbiters_next_2_5_sva | or_tmp_496;
  assign mux_405_nl = MUX_s_1_2_2(mux_404_nl, or_792_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_406_nl = MUX_s_1_2_2(or_tmp_496, mux_405_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign nor_623_nl = ~(and_1118_cse | and_1119_cse | mux_406_nl);
  assign mux_407_nl = MUX_s_1_2_2(nor_622_nl, nor_623_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl,
      mux_407_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1) & not_tmp_449;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 & not_tmp_449;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 | mux_450_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 & (~ mux_450_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1) & and_dcpl_720;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 & and_dcpl_720;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]),
      {mux_tmp_415 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1,
      {mux_tmp_415 , not_tmp_449 , (~ mux_450_itm) , and_dcpl_720});
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl,
      mux_tmp_440);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_4,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_5,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_6,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = (pe_manager_base_weight_sva_mx2[14:4])
      + PEManager_15U_GetWeightAddr_else_acc_3_1;
  assign PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1[10:0];
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_mx0w0
      = Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1);
  assign nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_3_mux_mx0w1
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1,
      operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1);
  assign nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_5_mux_mx0w3
      = MUX_s_1_2_2((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]),
      operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1) & and_dcpl_723;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 & and_dcpl_723;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_5_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_mx0w0,
      nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_3_mux_mx0w1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]),
      nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_5_mux_mx0w3,
      {weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp
      , and_dcpl_722 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      , and_dcpl_724});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1,
      {weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp
      , and_dcpl_722 , and_dcpl_723 , and_dcpl_724});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_tmp,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp
      = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_tmp
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp
      = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1 | (weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 | (weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1 | (weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1 | (weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 | (weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]));
  assign operator_7_false_1_operator_7_false_1_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 | (weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]));
  assign weight_read_addrs_0_3_0_lpi_1_dfm_4 = MUX_v_4_2_2(4'b0000, pe_manager_base_weight_sva_mx1_3_0,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_4_false_acc_sdt_sva_1 = conv_u2s_4_5(pe_config_num_manager_sva)
      + 5'b11111;
  assign operator_4_false_acc_sdt_sva_1 = nl_operator_4_false_acc_sdt_sva_1[4:0];
  assign while_and_1266_cse_1 = (~ while_if_and_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_if_and_tmp_1 = PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      = ~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl = start_PopNB_mioi_data_rsc_z_mxwt
      & pe_config_is_valid_sva & start_PopNB_mioi_return_rsc_z_mxwt;
  assign PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl = pe_config_is_zero_first_sva
      & pe_manager_zero_active_sva;
  assign PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl = ~(pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign PECore_UpdateFSM_switch_lp_mux1h_14_nl = MUX1HOT_s_1_4_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl,
      PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl, pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1,
      PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl, {PECore_UpdateFSM_switch_lp_and_7_itm_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_2_1 , PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_5_1});
  assign PECore_UpdateFSM_next_state_0_lpi_1_dfm_4 = PECore_UpdateFSM_switch_lp_mux1h_14_nl
      & PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  assign pe_config_UpdateManagerCounter_if_if_unequal_tmp = pe_config_output_counter_sva
      != (operator_8_false_acc_sdt_sva_1[7:0]);
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      = ~(pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]));
  assign input_write_req_valid_lpi_1_dfm_5 = PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      & PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1 = ~(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_144_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_111_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[127:120]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_144_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_159_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_127_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:120]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_159_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112_sva_1
      = MUX_v_8_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_111_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_127_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_150_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_102_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[55:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_150_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_165_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_118_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[55:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_165_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_sva_1
      = MUX_v_8_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_102_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_118_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_151_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_105_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[79:72]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_151_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_166_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_121_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[79:72]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_166_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_sva_1
      = MUX_v_8_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_105_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_121_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_152_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_104_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[71:64]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_152_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_167_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_120_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[71:64]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_167_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_sva_1
      = MUX_v_8_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_104_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_120_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420});
  assign while_and_40_tmp = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0,
      or_dcpl_295);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4, nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0,
      or_dcpl_295);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5, nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0,
      or_dcpl_295);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6, nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0,
      or_dcpl_295);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0,
      or_dcpl_295);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0,
      or_dcpl_295);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0,
      or_dcpl_295);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0,
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0,
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0,
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1 = and_319_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  assign nl_operator_16_false_acc_sdt_sva_1 = conv_u2s_8_9(pe_manager_num_input_sva)
      + 9'b111111111;
  assign operator_16_false_acc_sdt_sva_1 = nl_operator_16_false_acc_sdt_sva_1[8:0];
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1 = ~((state_mux_1_cse!=2'b00)
      | state_0_sva_mx1);
  assign PECore_UpdateFSM_switch_lp_and_2_tmp_1 = pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
      & PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
  assign PECore_UpdateFSM_switch_lp_nor_tmp_1 = ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_6 | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1
      | PECore_RunScale_PECore_RunScale_if_and_1_svs_1 | PECore_PushOutput_PECore_PushOutput_if_and_svs_1);
  assign PECore_UpdateFSM_switch_lp_not_31_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign act_port_reg_data_16_0_sva_dfm_3 = MUX_v_17_2_2(17'b00000000000000000, act_port_reg_data_16_0_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_31_nl);
  assign PECore_UpdateFSM_switch_lp_not_32_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign act_port_reg_data_176_160_sva_dfm_3 = MUX_v_17_2_2(17'b00000000000000000,
      act_port_reg_data_176_160_sva_dfm_1_1, PECore_UpdateFSM_switch_lp_not_32_nl);
  assign PECore_UpdateFSM_switch_lp_not_33_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign act_port_reg_data_208_192_sva_dfm_3 = MUX_v_17_2_2(17'b00000000000000000,
      act_port_reg_data_208_192_sva_dfm_1_1, PECore_UpdateFSM_switch_lp_not_33_nl);
  assign PECore_UpdateFSM_switch_lp_not_30_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign act_port_reg_data_240_224_sva_dfm_3 = MUX_v_17_2_2(17'b00000000000000000,
      act_port_reg_data_240_224_sva_dfm_1_1, PECore_UpdateFSM_switch_lp_not_30_nl);
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp
      = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2) | reg_rva_in_reg_rw_sva_2_cse
      | (~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp!=8'b00000000))) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7])));
  assign PECore_DecodeAxiWrite_switch_lp_or_5_cse_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  assign rva_out_reg_data_63_sva_dfm_7 = PECore_PushAxiRsp_mux_23_itm_1 & rva_in_reg_rw_sva_5;
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_1_0_sva_1 = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]!=2'b00));
  assign input_mem_banks_write_if_for_if_and_stg_1_1_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b01);
  assign input_mem_banks_write_if_for_if_and_stg_1_2_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b10);
  assign input_mem_banks_write_if_for_if_and_stg_1_3_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b11);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign nl_PEManager_15U_GetInputAddr_acc_nl = input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt
      + (pe_manager_base_input_sva[7:0]);
  assign PEManager_15U_GetInputAddr_acc_nl = nl_PEManager_15U_GetInputAddr_acc_nl[7:0];
  assign input_write_addrs_lpi_1_dfm_2 = PEManager_15U_GetInputAddr_acc_nl & ({{7{PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1}},
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1})
      & ({{7{PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1}}, PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1});
  assign input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1 = ~((input_write_addrs_lpi_1_dfm_2[1:0]!=2'b00));
  assign input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b01);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b10);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b11);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2
      | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_4 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0011);
  assign PECore_DecodeAxiRead_switch_lp_nor_13_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_not_185 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 =
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:1]!=15'b000000000000000));
  assign PECore_PushAxiRsp_if_asn_79 = (~ rva_in_reg_rw_sva_10) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_81 = rva_in_reg_rw_sva_10 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_83 = input_read_req_valid_lpi_1_dfm_1_10 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign weight_mem_run_3_for_5_asn_447 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_449 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_451 = (weight_read_addrs_7_lpi_1_dfm_3_2_0[2])
      & nor_681_cse & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_453 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_455 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_457 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_459 = (weight_read_addrs_5_lpi_1_dfm_3_2_0[2])
      & nor_690_cse & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_412 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_420 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign while_and_39_cse = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign PECore_PushAxiRsp_if_asn_87 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign PECore_PushAxiRsp_if_asn_89 = (~ rva_in_reg_rw_sva_5) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign PECore_PushAxiRsp_if_asn_91 = rva_in_reg_rw_sva_5 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign while_asn_1039 = rva_in_reg_rw_sva_5 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_1
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_44_itm_1
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_152 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_156 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_2
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_2
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign Arbiter_8U_Roundrobin_pick_1_mux_589_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1443_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_589_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_590_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1442_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_590_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_591_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1441_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_591_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_592_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1440_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_592_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_593_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1439_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_593_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_594_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1438_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_594_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1437_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1430_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_601_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1429_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_601_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_602_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1428_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_602_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_33_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_603_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1427_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_603_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_604_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1426_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_604_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_605_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1425_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_605_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_606_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1424_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_606_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_607_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1422_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_607_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_609_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1420_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_609_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_611_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1418_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_611_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_612_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1417_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_612_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1416_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_613_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1415_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_613_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_20_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_614_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1414_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_614_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_19_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_615_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1413_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_615_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_18_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_616_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1412_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_616_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_17_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_618_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1410_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_618_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_15_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1409_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_619_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1408_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_619_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_622_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1405_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_622_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_dcpl_2 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7
      | rva_in_reg_rw_sva_9);
  assign and_dcpl_4 = while_stage_0_11 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
  assign and_dcpl_5 = and_dcpl_4 & (~ rva_in_reg_rw_sva_st_1_9);
  assign and_dcpl_24 = while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9);
  assign and_dcpl_29 = while_stage_0_9 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  assign and_dcpl_30 = while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign and_dcpl_33 = while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_5_nl = (~ weight_mem_run_3_for_weight_mem_run_3_for_and_1_tmp) | (~ while_stage_0_5)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign or_4_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_run_3_for_land_2_lpi_1_dfm_1);
  assign mux_tmp = MUX_s_1_2_2(or_5_nl, or_4_nl, while_stage_0_6);
  assign nand_32_cse = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & rva_in_reg_rw_sva_st_1_5);
  assign or_11_nl = (~ while_stage_0_6) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_run_3_for_land_1_lpi_1_dfm_2);
  assign mux_3_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_2, (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign nand_nl = ~(while_stage_0_6 & mux_3_nl);
  assign mux_tmp_4 = MUX_s_1_2_2(or_11_nl, nand_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign and_dcpl_41 = while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign not_tmp_29 = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_run_3_for_land_1_lpi_1_dfm_2));
  assign or_13_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_1_lpi_1_dfm_2;
  assign mux_6_itm = MUX_s_1_2_2(not_tmp_29, or_13_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign and_dcpl_48 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign or_tmp_7 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_run_3_for_land_6_lpi_1_dfm_1);
  assign or_tmp_14 = Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp;
  assign and_782_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  assign and_784_cse = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign and_783_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  assign or_tmp_19 = and_782_cse | and_783_cse | and_784_cse;
  assign or_tmp_26 = Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp;
  assign and_785_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  assign and_786_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  assign and_787_cse = weight_mem_read_arbxbar_arbiters_next_6_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign or_tmp_32 = and_785_cse | and_786_cse | and_787_cse;
  assign and_dcpl_83 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_dcpl_90 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_92 = (((Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)
      | or_tmp_26) & and_dcpl_90;
  assign and_dcpl_94 = (((Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 |
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1)
      | or_tmp_14) & and_dcpl_90;
  assign or_79_cse = and_804_cse | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp;
  assign and_dcpl_96 = or_79_cse & and_dcpl_90;
  assign or_dcpl_40 = Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp;
  assign and_dcpl_98 = (and_803_cse | or_dcpl_40) & and_dcpl_90;
  assign and_dcpl_100 = (and_769_cse | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1)
      & and_dcpl_90;
  assign or_100_cse = and_774_cse | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  assign and_dcpl_102 = or_100_cse & and_dcpl_90;
  assign and_dcpl_104 = (and_802_cse | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1)
      & and_dcpl_90;
  assign and_dcpl_106 = (and_801_cse | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1)
      & and_dcpl_90;
  assign or_dcpl_75 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4);
  assign nor_404_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]));
  assign and_113_cse = (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) |
      (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]))) & (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]))) & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]))) & nor_404_cse;
  assign nor_405_cse = ~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]));
  assign and_120_cse = nor_405_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]))) & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])));
  assign nor_412_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]));
  assign nor_409_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]));
  assign nor_410_cse = ~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]));
  assign and_127_cse = nor_409_cse & nor_410_cse & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]))) & nor_412_cse;
  assign nor_413_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]));
  assign and_134_cse = nor_413_cse & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4])));
  assign and_141_cse = (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]) |
      (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])));
  assign or_dcpl_80 = and_141_cse | or_dcpl_75;
  assign and_148_cse = (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]) |
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])));
  assign nor_428_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]));
  assign nor_427_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]));
  assign and_162_cse = (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) |
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])));
  assign and_dcpl_163 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign and_dcpl_164 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]));
  assign and_dcpl_165 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign and_dcpl_166 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]));
  assign and_dcpl_167 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign and_dcpl_168 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign and_dcpl_169 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign and_dcpl_170 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign and_dcpl_172 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_180 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign and_dcpl_189 = and_dcpl_172 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]);
  assign and_dcpl_190 = and_dcpl_172 & and_dcpl_164;
  assign and_dcpl_192 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_193 = and_dcpl_166 & and_dcpl_172;
  assign and_dcpl_195 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_196 = and_dcpl_167 & and_dcpl_172;
  assign and_dcpl_197 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign and_dcpl_198 = and_dcpl_197 & while_stage_0_4;
  assign and_dcpl_199 = and_dcpl_168 & and_dcpl_172;
  assign and_dcpl_200 = and_dcpl_172 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]);
  assign and_dcpl_201 = and_dcpl_172 & and_dcpl_165;
  assign and_dcpl_202 = and_dcpl_172 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]);
  assign and_dcpl_203 = and_dcpl_172 & and_dcpl_163;
  assign and_dcpl_205 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_206 = and_dcpl_169 & and_dcpl_172;
  assign and_dcpl_208 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_209 = and_dcpl_170 & and_dcpl_172;
  assign and_dcpl_212 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign and_dcpl_216 = (state_2_1_sva==2'b01) & (~ state_0_sva) & and_666_cse;
  assign nor_433_nl = ~((state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt));
  assign or_193_nl = state_0_sva | (state_2_1_sva[1]);
  assign mux_28_nl = MUX_s_1_2_2(nor_433_nl, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_193_nl);
  assign and_dcpl_219 = mux_28_nl & (~(PECore_RunFSM_switch_lp_nor_tmp_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign and_dcpl_220 = rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign or_dcpl_151 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]!=2'b01);
  assign and_dcpl_223 = reg_rva_in_PopNB_mioi_iswt0_cse & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_226 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01);
  assign and_dcpl_227 = and_dcpl_226 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]))
      & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign and_dcpl_228 = and_dcpl_227 & and_dcpl_223 & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign and_dcpl_230 = and_dcpl_227 & and_dcpl_223 & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_160 = (~ while_stage_0_10) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  assign mux_30_nl = MUX_s_1_2_2((~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2])),
      (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign or_209_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])
      | (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_tmp_31 = MUX_s_1_2_2(mux_30_nl, or_209_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign or_tmp_47 = rva_in_reg_rw_sva_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1
      | rva_in_reg_rw_sva_st_1_4;
  assign nor_436_cse = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]!=2'b00));
  assign and_dcpl_260 = PECore_RunFSM_switch_lp_equal_tmp_1_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_789_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  assign or_tmp_75 = (~(and_789_cse | (~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]))
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_15_tmp)) |
      (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign or_tmp_87 = (~(and_1114_cse | (~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]))
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp)) |
      (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign nor_tmp_29 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  assign and_795_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  assign and_792_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  assign and_794_cse = weight_mem_read_arbxbar_arbiters_next_1_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign and_793_cse = weight_mem_read_arbxbar_arbiters_next_1_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign or_268_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])) | (~
      weight_mem_read_arbxbar_arbiters_next_1_4_sva) | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  assign mux_81_nl = MUX_s_1_2_2(or_268_nl, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      and_792_cse);
  assign mux_82_nl = MUX_s_1_2_2(mux_81_nl, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      and_793_cse);
  assign mux_83_nl = MUX_s_1_2_2(mux_82_nl, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      and_794_cse);
  assign mux_tmp_84 = MUX_s_1_2_2(mux_83_nl, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      and_795_cse);
  assign or_tmp_104 = (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])))
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign and_dcpl_277 = while_stage_0_8 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6);
  assign and_dcpl_279 = while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6;
  assign and_dcpl_280 = while_stage_0_10 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  assign and_dcpl_281 = and_dcpl_220 & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_295 = and_dcpl_280 & (~ rva_in_reg_rw_sva_st_1_8);
  assign and_dcpl_308 = and_dcpl_295 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6
      | input_read_req_valid_lpi_1_dfm_1_8 | rva_in_reg_rw_sva_8));
  assign and_dcpl_314 = (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8) & PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
  assign and_dcpl_321 = and_dcpl_226 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]));
  assign and_dcpl_346 = and_dcpl_29 & (~ rva_in_reg_rw_sva_st_1_7);
  assign and_dcpl_351 = while_stage_0_9 & (~ rva_in_reg_rw_sva_7);
  assign and_dcpl_359 = and_dcpl_351 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & (~(rva_in_reg_rw_sva_st_1_7 | input_read_req_valid_lpi_1_dfm_1_7 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5));
  assign and_dcpl_370 = and_dcpl_279 & (~ rva_in_reg_rw_sva_st_1_6);
  assign and_dcpl_373 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4
      | rva_in_reg_rw_sva_6 | input_read_req_valid_lpi_1_dfm_1_6);
  assign and_dcpl_374 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
      & (~ rva_in_reg_rw_sva_st_1_6);
  assign and_dcpl_399 = ~(rva_in_reg_rw_sva_st_1_5 | rva_in_reg_rw_sva_5 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_dcpl_403 = and_dcpl_41 & (~ rva_in_reg_rw_sva_st_1_5);
  assign nand_40_cse = ~(while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_tmp_115 = (~ while_stage_0_5) | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | rva_in_reg_rw_sva_3;
  assign and_dcpl_433 = (~ rva_in_reg_rw_sva_3) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_dcpl_434 = (~ input_read_req_valid_lpi_1_dfm_1_3) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2;
  assign and_dcpl_435 = ~(pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1);
  assign or_dcpl_201 = crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp | (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp);
  assign and_dcpl_458 = or_dcpl_201 & (~(reg_rva_in_reg_rw_sva_2_cse | input_read_req_valid_lpi_1_dfm_1_2));
  assign and_dcpl_479 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | input_read_req_valid_lpi_1_dfm_1_1);
  assign and_dcpl_480 = and_dcpl_479 & and_dcpl_212;
  assign mux_tmp_110 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1!=4'b0100));
  assign and_dcpl_488 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1);
  assign nand_41_cse = ~(PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]));
  assign and_dcpl_524 = PECore_RunMac_PECore_RunMac_if_and_svs_st_6 & while_stage_0_8
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6);
  assign and_dcpl_528 = while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
  assign and_dcpl_534 = and_dcpl_83 & (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign or_332_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1;
  assign mux_111_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      or_332_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_tmp_1 = while_stage_0_6 & mux_111_nl;
  assign and_dcpl_537 = (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign or_336_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1;
  assign mux_113_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      or_336_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_tmp_2 = while_stage_0_6 & mux_113_nl;
  assign or_341_nl = Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse;
  assign mux_tmp_115 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1,
      or_341_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_340_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign mux_116_nl = MUX_s_1_2_2(mux_tmp_115, or_340_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_3 = while_stage_0_5 & mux_116_nl;
  assign and_547_nl = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 & (Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse);
  assign or_347_nl = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1;
  assign mux_119_nl = MUX_s_1_2_2(and_547_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1,
      or_347_nl);
  assign or_tmp_136 = Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 | mux_119_nl;
  assign or_346_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign mux_120_nl = MUX_s_1_2_2(or_tmp_136, or_346_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_5 = while_stage_0_5 & mux_120_nl;
  assign and_dcpl_545 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign or_352_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign mux_123_nl = MUX_s_1_2_2(or_100_cse, or_352_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_7 = while_stage_0_5 & mux_123_nl;
  assign or_360_nl = Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6;
  assign mux_tmp_126 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1,
      or_360_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_359_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_3 | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign mux_127_nl = MUX_s_1_2_2(mux_tmp_126, or_359_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_8 = while_stage_0_5 & mux_127_nl;
  assign or_363_nl = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  assign mux_tmp_130 = MUX_s_1_2_2(or_dcpl_40, or_363_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign mux_tmp_131 = MUX_s_1_2_2(mux_tmp_130, PECore_RunMac_PECore_RunMac_if_and_svs_st_3,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_562_nl = while_stage_0_5 & mux_tmp_131;
  assign and_561_nl = while_stage_0_5 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | mux_tmp_130);
  assign mux_tmp_132 = MUX_s_1_2_2(and_562_nl, and_561_nl, PECore_UpdateFSM_switch_lp_equal_tmp_2_3);
  assign or_370_nl = PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 | PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign mux_135_nl = MUX_s_1_2_2(or_79_cse, or_370_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_11 = while_stage_0_5 & mux_135_nl;
  assign and_dcpl_561 = fsm_output & (~ weight_mem_run_3_for_land_5_lpi_1_dfm_3);
  assign and_dcpl_562 = fsm_output & (~ weight_mem_run_3_for_land_3_lpi_1_dfm_3);
  assign or_dcpl_220 = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_9) | PECore_RunMac_PECore_RunMac_if_and_svs_st_9;
  assign or_dcpl_221 = (~ while_stage_0_8) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6;
  assign or_dcpl_227 = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign and_dcpl_578 = or_dcpl_227 & weight_mem_run_3_for_land_1_lpi_1_dfm_3 & (~
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_dcpl_580 = or_dcpl_227 & (~(weight_mem_run_3_for_land_1_lpi_1_dfm_3
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5));
  assign and_dcpl_581 = or_dcpl_227 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign and_dcpl_583 = and_dcpl_48 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign or_dcpl_231 = (~ while_stage_0_7) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign or_dcpl_233 = or_dcpl_231 | (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign and_dcpl_600 = and_dcpl_90 & (~ while_stage_0_4);
  assign or_dcpl_236 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ while_stage_0_5);
  assign and_dcpl_643 = (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]) |
      (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]))) & nor_427_cse & nor_428_cse;
  assign or_dcpl_237 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ while_stage_0_3);
  assign or_dcpl_249 = or_dcpl_151 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]);
  assign or_dcpl_256 = nand_88_cse | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_257 = (~ while_stage_0_12) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10;
  assign and_dcpl_655 = or_dcpl_227 & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign and_dcpl_656 = or_dcpl_227 & (~ weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign and_dcpl_657 = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]==2'b10);
  assign and_dcpl_659 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign and_dcpl_660 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]));
  assign and_dcpl_661 = and_dcpl_660 & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign and_dcpl_662 = and_dcpl_660 & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]));
  assign and_dcpl_663 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign and_dcpl_670 = ~(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_dcpl_284 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | nand_41_cse;
  assign or_dcpl_287 = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_8) | PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
  assign or_dcpl_291 = (~(while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6))
      | rva_in_reg_rw_sva_6;
  assign nor_tmp_53 = weight_mem_read_arbxbar_arbiters_next_7_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign or_tmp_172 = and_782_cse | nor_tmp_53;
  assign or_466_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign mux_tmp_160 = MUX_s_1_2_2(or_tmp_172, or_466_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign nor_tmp_55 = Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign and_813_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) & Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1;
  assign or_469_cse = and_813_cse | nor_tmp_55;
  assign mux_tmp_161 = MUX_s_1_2_2(or_tmp_172, or_469_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign mux_164_nl = MUX_s_1_2_2(mux_tmp_161, mux_tmp_160, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_165_nl = MUX_s_1_2_2(or_tmp_172, mux_164_nl, while_stage_0_5);
  assign or_471_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | or_tmp_172;
  assign or_470_nl = Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 | mux_tmp_161;
  assign or_468_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | mux_tmp_160;
  assign mux_162_nl = MUX_s_1_2_2(or_470_nl, or_468_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_163_nl = MUX_s_1_2_2(or_471_nl, mux_162_nl, while_stage_0_5);
  assign mux_tmp_166 = MUX_s_1_2_2(mux_165_nl, mux_163_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign nand_tmp_7 = ~(weight_mem_read_arbxbar_arbiters_next_7_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      & (~ or_tmp_172));
  assign and_817_cse = weight_mem_read_arbxbar_arbiters_next_7_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign mux_170_nl = MUX_s_1_2_2(nand_tmp_7, or_tmp_172, and_817_cse);
  assign mux_168_nl = MUX_s_1_2_2(nand_tmp_7, or_tmp_172, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign or_475_nl = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign mux_167_nl = MUX_s_1_2_2(nand_tmp_7, or_tmp_172, or_475_nl);
  assign mux_169_nl = MUX_s_1_2_2(mux_168_nl, mux_167_nl, weight_mem_read_arbxbar_arbiters_next_7_3_sva);
  assign mux_171_nl = MUX_s_1_2_2(mux_170_nl, mux_169_nl, weight_mem_read_arbxbar_arbiters_next_7_2_sva);
  assign mux_tmp_172 = MUX_s_1_2_2(mux_171_nl, or_tmp_172, and_797_cse);
  assign and_824_cse = Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign and_826_cse = Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign and_825_cse = Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign nor_551_nl = ~(and_784_cse | mux_tmp_172);
  assign nand_8_nl = ~(Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      & (~ or_469_cse));
  assign mux_174_nl = MUX_s_1_2_2(nand_8_nl, or_469_cse, and_824_cse);
  assign mux_175_nl = MUX_s_1_2_2(mux_174_nl, or_469_cse, and_825_cse);
  assign mux_176_nl = MUX_s_1_2_2(mux_175_nl, or_469_cse, and_826_cse);
  assign mux_177_nl = MUX_s_1_2_2(mux_tmp_172, mux_176_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign nor_552_nl = ~((Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]))
      | mux_177_nl);
  assign or_473_nl = (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])))
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign mux_173_nl = MUX_s_1_2_2(mux_tmp_172, or_473_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign nor_553_nl = ~(and_784_cse | mux_173_nl);
  assign mux_178_nl = MUX_s_1_2_2(nor_552_nl, nor_553_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign not_tmp_404 = MUX_s_1_2_2(nor_551_nl, mux_178_nl, while_stage_0_5);
  assign or_tmp_187 = and_783_cse | and_817_cse | nor_tmp_53;
  assign or_tmp_190 = and_797_cse | and_798_cse | and_782_cse | or_tmp_187;
  assign or_480_nl = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign mux_tmp_180 = MUX_s_1_2_2(or_tmp_190, or_480_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign and_833_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) & Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1;
  assign or_tmp_193 = and_833_cse | and_824_cse | nor_tmp_55;
  assign or_491_nl = and_826_cse | and_825_cse | and_813_cse | or_tmp_193;
  assign mux_tmp_181 = MUX_s_1_2_2(or_tmp_190, or_491_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_493_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | or_tmp_190;
  assign or_492_nl = Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 | mux_tmp_181;
  assign or_486_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | mux_tmp_180;
  assign mux_182_nl = MUX_s_1_2_2(or_492_nl, or_486_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_183 = MUX_s_1_2_2(or_493_nl, mux_182_nl, while_stage_0_5);
  assign mux_184_nl = MUX_s_1_2_2(mux_tmp_181, mux_tmp_180, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_185 = MUX_s_1_2_2(or_tmp_190, mux_184_nl, while_stage_0_5);
  assign or_497_nl = and_783_cse | and_817_cse | weight_mem_read_arbxbar_arbiters_next_7_6_sva
      | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]));
  assign or_494_nl = weight_mem_read_arbxbar_arbiters_next_7_5_sva | or_tmp_187;
  assign mux_186_nl = MUX_s_1_2_2(or_497_nl, or_494_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign or_tmp_204 = and_797_cse | and_798_cse | mux_186_nl;
  assign or_504_nl = and_833_cse | and_824_cse | Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1
      | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]));
  assign or_501_nl = Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 | or_tmp_193;
  assign mux_187_nl = MUX_s_1_2_2(or_504_nl, or_501_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign or_506_nl = and_826_cse | and_825_cse | mux_187_nl;
  assign mux_188_nl = MUX_s_1_2_2(or_tmp_204, or_506_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_500_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7])
      | or_tmp_204;
  assign mux_189_nl = MUX_s_1_2_2(mux_188_nl, or_500_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_190_nl = MUX_s_1_2_2(or_tmp_204, mux_189_nl, while_stage_0_5);
  assign mux_191_nl = MUX_s_1_2_2(mux_190_nl, mux_tmp_185, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign mux_192_itm = MUX_s_1_2_2(mux_191_nl, mux_tmp_183, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign or_tmp_212 = and_783_cse | and_817_cse;
  assign or_512_nl = weight_mem_read_arbxbar_arbiters_next_7_3_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]));
  assign or_511_nl = weight_mem_read_arbxbar_arbiters_next_7_4_sva | and_817_cse;
  assign mux_193_nl = MUX_s_1_2_2(or_512_nl, or_511_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign or_510_nl = weight_mem_read_arbxbar_arbiters_next_7_2_sva | or_tmp_212;
  assign mux_194_nl = MUX_s_1_2_2(mux_193_nl, or_510_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign or_509_nl = weight_mem_read_arbxbar_arbiters_next_7_1_sva | and_798_cse
      | or_tmp_212;
  assign mux_tmp_195 = MUX_s_1_2_2(mux_194_nl, or_509_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign or_tmp_219 = and_833_cse | and_824_cse;
  assign or_519_nl = Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]));
  assign or_518_nl = Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 | and_824_cse;
  assign mux_196_nl = MUX_s_1_2_2(or_519_nl, or_518_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign or_517_nl = Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 | or_tmp_219;
  assign mux_197_nl = MUX_s_1_2_2(mux_196_nl, or_517_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign or_516_nl = Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 | and_825_cse | or_tmp_219;
  assign mux_198_nl = MUX_s_1_2_2(mux_197_nl, or_516_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign mux_199_nl = MUX_s_1_2_2(mux_tmp_195, mux_198_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_513_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7])
      | mux_tmp_195;
  assign mux_200_nl = MUX_s_1_2_2(mux_199_nl, or_513_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_201_nl = MUX_s_1_2_2(mux_tmp_195, mux_200_nl, while_stage_0_5);
  assign and_dcpl_698 = (~ mux_201_nl) & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]))) & nor_404_cse;
  assign and_853_cse = while_mux_1437_tmp & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_tmp_225 = ((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & while_mux_1439_tmp)
      | and_853_cse;
  assign or_tmp_227 = and_785_cse | (Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]));
  assign mux_204_nl = MUX_s_1_2_2(or_tmp_227, or_tmp_225, while_stage_0_5);
  assign or_523_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | or_tmp_227;
  assign or_521_nl = while_mux_1438_tmp | or_tmp_225;
  assign mux_203_nl = MUX_s_1_2_2(or_523_nl, or_521_nl, while_stage_0_5);
  assign mux_tmp_205 = MUX_s_1_2_2(mux_204_nl, mux_203_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign and_859_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & while_mux_1442_tmp;
  assign and_857_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]) & while_mux_1443_tmp;
  assign and_858_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & while_mux_1441_tmp;
  assign nand_9_nl = ~(while_mux_1440_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      & (~ or_tmp_225));
  assign mux_206_nl = MUX_s_1_2_2(nand_9_nl, or_tmp_225, and_857_cse);
  assign mux_207_nl = MUX_s_1_2_2(mux_206_nl, or_tmp_225, and_858_cse);
  assign mux_tmp_208 = MUX_s_1_2_2(mux_207_nl, or_tmp_225, and_859_cse);
  assign and_862_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  assign nand_10_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      & (~ or_tmp_227));
  assign mux_209_nl = MUX_s_1_2_2(nand_10_nl, or_tmp_227, and_799_cse);
  assign mux_210_nl = MUX_s_1_2_2(mux_209_nl, or_tmp_227, and_862_cse);
  assign mux_tmp_211 = MUX_s_1_2_2(mux_210_nl, or_tmp_227, and_800_cse);
  assign mux_213_nl = MUX_s_1_2_2(mux_tmp_211, mux_tmp_208, while_stage_0_5);
  assign or_525_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | mux_tmp_211;
  assign or_524_nl = while_mux_1438_tmp | mux_tmp_208;
  assign mux_212_nl = MUX_s_1_2_2(or_525_nl, or_524_nl, while_stage_0_5);
  assign mux_214_itm = MUX_s_1_2_2(mux_213_nl, mux_212_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign nor_tmp_109 = while_mux_1438_tmp & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign or_tmp_232 = and_853_cse | nor_tmp_109;
  assign and_867_cse = while_mux_1440_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign or_530_nl = while_mux_1438_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign or_529_nl = while_mux_1437_tmp | nor_tmp_109;
  assign mux_215_nl = MUX_s_1_2_2(or_530_nl, or_529_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_216_nl = MUX_s_1_2_2(mux_215_nl, or_tmp_232, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_528_nl = while_mux_1439_tmp | or_tmp_232;
  assign mux_217_nl = MUX_s_1_2_2(mux_216_nl, or_528_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_237 = and_859_cse | and_867_cse | mux_217_nl;
  assign or_tmp_240 = and_786_cse | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  assign mux_tmp_218 = MUX_s_1_2_2(and_786_cse, or_tmp_240, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_537_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign mux_219_nl = MUX_s_1_2_2(or_537_nl, or_tmp_240, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_220_nl = MUX_s_1_2_2(mux_219_nl, mux_tmp_218, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_536_nl = weight_mem_read_arbxbar_arbiters_next_6_5_sva | mux_tmp_218;
  assign mux_221_nl = MUX_s_1_2_2(mux_220_nl, or_536_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_244 = and_800_cse | and_787_cse | mux_221_nl;
  assign mux_226_nl = MUX_s_1_2_2(or_tmp_244, or_tmp_237, while_stage_0_5);
  assign or_544_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | or_tmp_244;
  assign or_543_nl = while_mux_1441_tmp | or_tmp_237;
  assign mux_225_nl = MUX_s_1_2_2(or_544_nl, or_543_nl, while_stage_0_5);
  assign mux_227_nl = MUX_s_1_2_2(mux_226_nl, mux_225_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign or_542_nl = weight_mem_read_arbxbar_arbiters_next_6_1_sva | or_tmp_244;
  assign or_541_nl = while_mux_1443_tmp | or_tmp_237;
  assign mux_223_nl = MUX_s_1_2_2(or_542_nl, or_541_nl, while_stage_0_5);
  assign or_540_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | or_tmp_244;
  assign or_533_nl = while_mux_1441_tmp | while_mux_1443_tmp | or_tmp_237;
  assign mux_222_nl = MUX_s_1_2_2(or_540_nl, or_533_nl, while_stage_0_5);
  assign mux_224_nl = MUX_s_1_2_2(mux_223_nl, mux_222_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_228_itm = MUX_s_1_2_2(mux_227_nl, mux_224_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_tmp_250 = and_857_cse | and_867_cse;
  assign or_tmp_256 = and_799_cse | and_787_cse;
  assign nor_555_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])));
  assign nor_556_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_1_sva | and_787_cse);
  assign mux_232_nl = MUX_s_1_2_2(nor_555_nl, nor_556_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign nor_557_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_3_sva | or_tmp_256);
  assign mux_233_nl = MUX_s_1_2_2(mux_232_nl, nor_557_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nor_558_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_2_sva | and_862_cse
      | or_tmp_256);
  assign mux_234_nl = MUX_s_1_2_2(mux_233_nl, nor_558_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign nor_559_nl = ~(while_mux_1440_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])));
  assign nor_560_nl = ~(while_mux_1443_tmp | and_867_cse);
  assign mux_229_nl = MUX_s_1_2_2(nor_559_nl, nor_560_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign nor_561_nl = ~(while_mux_1441_tmp | or_tmp_250);
  assign mux_230_nl = MUX_s_1_2_2(mux_229_nl, nor_561_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nor_562_nl = ~(while_mux_1442_tmp | and_858_cse | or_tmp_250);
  assign mux_231_nl = MUX_s_1_2_2(mux_230_nl, nor_562_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign mux_235_nl = MUX_s_1_2_2(mux_234_nl, mux_231_nl, while_stage_0_5);
  assign and_dcpl_701 = mux_235_nl & nor_405_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])));
  assign or_tmp_265 = and_859_cse | and_858_cse | and_857_cse | and_867_cse | or_tmp_225;
  assign or_tmp_270 = and_800_cse | and_862_cse | and_799_cse | and_787_cse | or_tmp_227;
  assign and_887_cse = weight_mem_read_arbxbar_arbiters_next_5_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign and_886_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  assign or_tmp_273 = and_886_cse | and_887_cse;
  assign or_569_cse = and_1100_cse | and_1101_cse;
  assign mux_240_nl = MUX_s_1_2_2(or_tmp_273, or_569_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_567_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign mux_239_nl = MUX_s_1_2_2(or_tmp_273, or_567_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign mux_tmp_241 = MUX_s_1_2_2(mux_240_nl, mux_239_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_243_nl = MUX_s_1_2_2(or_tmp_273, mux_tmp_241, while_stage_0_5);
  assign or_571_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1
      | or_tmp_273;
  assign or_570_nl = while_mux_1430_tmp | mux_tmp_241;
  assign mux_242_nl = MUX_s_1_2_2(or_571_nl, or_570_nl, while_stage_0_5);
  assign mux_tmp_244 = MUX_s_1_2_2(mux_243_nl, mux_242_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign and_895_cse = weight_mem_read_arbxbar_arbiters_next_5_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign nand_11_nl = ~(weight_mem_read_arbxbar_arbiters_next_5_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      & (~ or_tmp_273));
  assign mux_248_cse = MUX_s_1_2_2(nand_11_nl, or_tmp_273, and_895_cse);
  assign mux_255_nl = MUX_s_1_2_2(mux_248_cse, or_tmp_273, and_1094_cse);
  assign mux_256_nl = MUX_s_1_2_2(mux_255_nl, or_tmp_273, and_1093_cse);
  assign nor_565_nl = ~(and_1092_cse | mux_256_nl);
  assign nand_12_nl = ~(Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      & (~ or_569_cse));
  assign mux_250_nl = MUX_s_1_2_2(nand_12_nl, or_569_cse, and_1098_cse);
  assign mux_251_nl = MUX_s_1_2_2(mux_248_cse, mux_250_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_576_nl = nor_410_cse | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign mux_249_nl = MUX_s_1_2_2(mux_248_cse, or_576_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign mux_252_nl = MUX_s_1_2_2(mux_251_nl, mux_249_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_253_nl = MUX_s_1_2_2(mux_252_nl, mux_tmp_241, and_1097_cse);
  assign mux_254_nl = MUX_s_1_2_2(mux_253_nl, mux_tmp_241, and_1096_cse);
  assign nor_566_nl = ~(and_1095_cse | mux_254_nl);
  assign not_tmp_417 = MUX_s_1_2_2(nor_565_nl, nor_566_nl, while_stage_0_5);
  assign and_906_cse = weight_mem_read_arbxbar_arbiters_next_5_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign or_tmp_287 = and_895_cse | and_906_cse | and_886_cse | and_887_cse;
  assign or_593_nl = weight_mem_read_arbxbar_arbiters_next_5_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]));
  assign or_592_nl = weight_mem_read_arbxbar_arbiters_next_5_5_sva | and_887_cse;
  assign mux_262_nl = MUX_s_1_2_2(or_593_nl, or_592_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign or_tmp_300 = and_895_cse | and_906_cse | mux_262_nl;
  assign mux_267_nl = MUX_s_1_2_2(or_tmp_300, or_tmp_287, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign nor_567_nl = ~(and_1093_cse | and_1094_cse | mux_267_nl);
  assign or_598_nl = Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]));
  assign or_597_nl = Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 | and_1101_cse;
  assign mux_263_nl = MUX_s_1_2_2(or_598_nl, or_597_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign or_600_nl = and_1098_cse | and_1099_cse | mux_263_nl;
  assign mux_264_nl = MUX_s_1_2_2(or_tmp_300, or_600_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_596_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5])
      | or_tmp_300;
  assign mux_265_nl = MUX_s_1_2_2(mux_264_nl, or_596_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_266_nl = MUX_s_1_2_2(mux_265_nl, mux_285_cse, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign nor_568_nl = ~(and_1096_cse | and_1097_cse | mux_266_nl);
  assign mux_268_nl = MUX_s_1_2_2(nor_567_nl, nor_568_nl, while_stage_0_5);
  assign nor_569_nl = ~(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1
      | and_1093_cse | and_1094_cse | or_tmp_287);
  assign nor_570_nl = ~(while_mux_1430_tmp | and_1096_cse | and_1097_cse | mux_285_cse);
  assign mux_261_nl = MUX_s_1_2_2(nor_569_nl, nor_570_nl, while_stage_0_5);
  assign not_tmp_419 = MUX_s_1_2_2(mux_268_nl, mux_261_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign or_tmp_311 = and_895_cse | and_906_cse;
  assign mux_tmp_270 = MUX_s_1_2_2(or_tmp_311, operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1,
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign or_611_nl = weight_mem_read_arbxbar_arbiters_next_5_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]));
  assign or_610_nl = weight_mem_read_arbxbar_arbiters_next_5_3_sva | and_906_cse;
  assign mux_tmp_271 = MUX_s_1_2_2(or_611_nl, or_610_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign or_613_nl = and_1098_cse | and_1099_cse;
  assign mux_tmp_274 = MUX_s_1_2_2(or_tmp_311, or_613_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_621_nl = weight_mem_read_arbxbar_arbiters_next_5_2_sva | or_tmp_311;
  assign mux_280_nl = MUX_s_1_2_2(mux_tmp_271, or_621_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign or_620_nl = weight_mem_read_arbxbar_arbiters_next_5_1_sva | and_1094_cse
      | or_tmp_311;
  assign mux_281_nl = MUX_s_1_2_2(mux_280_nl, or_620_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign or_618_nl = Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]));
  assign or_617_nl = Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 | and_1099_cse;
  assign mux_275_nl = MUX_s_1_2_2(or_618_nl, or_617_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign mux_276_nl = MUX_s_1_2_2(mux_tmp_271, mux_275_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_616_nl = Arbiter_8U_Roundrobin_pick_1_mux_428_mx1w1 | mux_tmp_274;
  assign mux_277_nl = MUX_s_1_2_2(mux_276_nl, or_616_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign or_615_nl = Arbiter_8U_Roundrobin_pick_1_mux_429_mx1w1 | ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5])
      & Arbiter_8U_Roundrobin_pick_1_mux_428_mx1w1) | mux_tmp_274;
  assign mux_278_nl = MUX_s_1_2_2(mux_277_nl, or_615_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign or_612_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5])
      | mux_tmp_271;
  assign or_609_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0
      | mux_tmp_270;
  assign mux_272_nl = MUX_s_1_2_2(or_612_nl, or_609_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign or_608_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0
      | ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0)
      | mux_tmp_270;
  assign mux_273_nl = MUX_s_1_2_2(mux_272_nl, or_608_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign mux_279_nl = MUX_s_1_2_2(mux_278_nl, mux_273_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_282_nl = MUX_s_1_2_2(mux_281_nl, mux_279_nl, while_stage_0_5);
  assign and_dcpl_703 = (~ mux_282_nl) & nor_409_cse & nor_412_cse;
  assign nor_tmp_189 = while_mux_1425_tmp & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign and_937_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1;
  assign and_939_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) & while_mux_1424_tmp;
  assign and_940_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]) & Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1;
  assign and_938_cse = weight_mem_read_arbxbar_arbiters_next_4_5_sva & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign and_936_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  assign or_639_cse = and_936_cse | and_937_cse | and_938_cse;
  assign or_636_nl = and_940_cse | nor_tmp_189;
  assign or_635_nl = and_937_cse | nor_tmp_189;
  assign mux_287_nl = MUX_s_1_2_2(or_636_nl, or_635_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_637_nl = and_939_cse | mux_287_nl;
  assign mux_tmp_288 = MUX_s_1_2_2(or_639_cse, or_637_nl, while_stage_0_5);
  assign or_tmp_345 = while_mux_1427_tmp | while_mux_1429_tmp;
  assign mux_289_cse = MUX_s_1_2_2(and_940_cse, and_937_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_347 = nor_tmp_189 | and_939_cse | mux_289_cse;
  assign and_947_cse = while_mux_1428_tmp & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign or_tmp_348 = weight_mem_read_arbxbar_arbiters_next_4_1_sva | weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  assign and_951_cse = weight_mem_read_arbxbar_arbiters_next_4_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign nand_14_nl = ~(weight_mem_read_arbxbar_arbiters_next_4_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])
      & (~ or_639_cse));
  assign mux_292_itm = MUX_s_1_2_2(nand_14_nl, or_639_cse, and_951_cse);
  assign nand_13_nl = ~(while_mux_1426_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])
      & (~ or_tmp_347));
  assign mux_290_itm = MUX_s_1_2_2(nand_13_nl, or_tmp_347, and_947_cse);
  assign mux_302_nl = MUX_s_1_2_2(mux_292_itm, mux_290_itm, while_stage_0_5);
  assign mux_300_nl = MUX_s_1_2_2(mux_292_itm, or_639_cse, weight_mem_read_arbxbar_arbiters_next_4_3_sva);
  assign mux_299_nl = MUX_s_1_2_2(mux_290_itm, or_tmp_347, while_mux_1427_tmp);
  assign mux_301_nl = MUX_s_1_2_2(mux_300_nl, mux_299_nl, while_stage_0_5);
  assign mux_303_nl = MUX_s_1_2_2(mux_302_nl, mux_301_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign mux_296_nl = MUX_s_1_2_2(mux_292_itm, or_639_cse, weight_mem_read_arbxbar_arbiters_next_4_1_sva);
  assign mux_295_nl = MUX_s_1_2_2(mux_290_itm, or_tmp_347, while_mux_1429_tmp);
  assign mux_297_nl = MUX_s_1_2_2(mux_296_nl, mux_295_nl, while_stage_0_5);
  assign mux_293_nl = MUX_s_1_2_2(mux_292_itm, or_639_cse, or_tmp_348);
  assign mux_291_nl = MUX_s_1_2_2(mux_290_itm, or_tmp_347, or_tmp_345);
  assign mux_294_nl = MUX_s_1_2_2(mux_293_nl, mux_291_nl, while_stage_0_5);
  assign mux_298_nl = MUX_s_1_2_2(mux_297_nl, mux_294_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign mux_304_itm = MUX_s_1_2_2(mux_303_nl, mux_298_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign mux_305_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_353 = nor_tmp_189 | and_939_cse | mux_305_nl;
  assign or_651_nl = while_mux_1424_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]));
  assign mux_306_nl = MUX_s_1_2_2(or_651_nl, and_939_cse, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]);
  assign or_650_nl = while_mux_1425_tmp | and_939_cse;
  assign mux_tmp_307 = MUX_s_1_2_2(mux_306_nl, or_650_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign mux_309_nl = MUX_s_1_2_2(mux_tmp_307, or_tmp_353, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign or_652_nl = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | mux_tmp_307;
  assign or_649_nl = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | or_tmp_353;
  assign mux_308_nl = MUX_s_1_2_2(or_652_nl, or_649_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign mux_310_nl = MUX_s_1_2_2(mux_309_nl, mux_308_nl, while_mux_1426_tmp);
  assign or_tmp_358 = and_947_cse | mux_310_nl;
  assign or_tmp_362 = and_938_cse | and_936_cse | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1;
  assign or_660_nl = weight_mem_read_arbxbar_arbiters_next_4_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]));
  assign mux_311_nl = MUX_s_1_2_2(or_660_nl, and_936_cse, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]);
  assign or_659_nl = weight_mem_read_arbxbar_arbiters_next_4_5_sva | and_936_cse;
  assign mux_tmp_312 = MUX_s_1_2_2(mux_311_nl, or_659_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign mux_314_nl = MUX_s_1_2_2(mux_tmp_312, or_tmp_362, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign or_661_nl = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | mux_tmp_312;
  assign or_658_nl = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | or_tmp_362;
  assign mux_313_nl = MUX_s_1_2_2(or_661_nl, or_658_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign mux_315_nl = MUX_s_1_2_2(mux_314_nl, mux_313_nl, weight_mem_read_arbxbar_arbiters_next_4_4_sva);
  assign or_tmp_367 = and_951_cse | mux_315_nl;
  assign mux_320_nl = MUX_s_1_2_2(or_tmp_367, or_tmp_358, while_stage_0_5);
  assign or_667_nl = weight_mem_read_arbxbar_arbiters_next_4_3_sva | or_tmp_367;
  assign or_666_nl = while_mux_1427_tmp | or_tmp_358;
  assign mux_319_nl = MUX_s_1_2_2(or_667_nl, or_666_nl, while_stage_0_5);
  assign mux_321_nl = MUX_s_1_2_2(mux_320_nl, mux_319_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign or_665_nl = weight_mem_read_arbxbar_arbiters_next_4_1_sva | or_tmp_367;
  assign or_664_nl = while_mux_1429_tmp | or_tmp_358;
  assign mux_317_nl = MUX_s_1_2_2(or_665_nl, or_664_nl, while_stage_0_5);
  assign or_663_nl = or_tmp_348 | or_tmp_367;
  assign or_654_nl = or_tmp_345 | or_tmp_358;
  assign mux_316_nl = MUX_s_1_2_2(or_663_nl, or_654_nl, while_stage_0_5);
  assign mux_318_nl = MUX_s_1_2_2(mux_317_nl, mux_316_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign mux_322_itm = MUX_s_1_2_2(mux_321_nl, mux_318_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign nor_tmp_214 = while_mux_1427_tmp & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign or_tmp_373 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]) & while_mux_1429_tmp)
      | nor_tmp_214;
  assign nor_tmp_217 = weight_mem_read_arbxbar_arbiters_next_4_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign or_tmp_379 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_1_sva)
      | nor_tmp_217;
  assign nor_571_nl = ~(weight_mem_read_arbxbar_arbiters_next_4_3_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])));
  assign nor_572_nl = ~(weight_mem_read_arbxbar_arbiters_next_4_1_sva | nor_tmp_217);
  assign mux_326_nl = MUX_s_1_2_2(nor_571_nl, nor_572_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign nor_573_nl = ~(weight_mem_read_arbxbar_arbiters_next_4_2_sva | or_tmp_379);
  assign mux_327_nl = MUX_s_1_2_2(mux_326_nl, nor_573_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign nor_574_nl = ~(weight_mem_read_arbxbar_arbiters_next_4_4_sva | and_951_cse
      | or_tmp_379);
  assign mux_328_nl = MUX_s_1_2_2(mux_327_nl, nor_574_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign nor_575_nl = ~(while_mux_1427_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])));
  assign nor_576_nl = ~(while_mux_1429_tmp | nor_tmp_214);
  assign mux_323_nl = MUX_s_1_2_2(nor_575_nl, nor_576_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign nor_577_nl = ~(while_mux_1428_tmp | or_tmp_373);
  assign mux_324_nl = MUX_s_1_2_2(mux_323_nl, nor_577_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign nor_578_nl = ~(while_mux_1426_tmp | and_947_cse | or_tmp_373);
  assign mux_325_nl = MUX_s_1_2_2(mux_324_nl, nor_578_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign mux_329_nl = MUX_s_1_2_2(mux_328_nl, mux_325_nl, while_stage_0_5);
  assign and_dcpl_706 = mux_329_nl & nor_413_cse & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4])));
  assign or_tmp_389 = and_947_cse | (while_mux_1426_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]))
      | nor_tmp_189 | and_939_cse | mux_289_cse;
  assign or_tmp_395 = and_951_cse | (weight_mem_read_arbxbar_arbiters_next_4_4_sva
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])) | and_938_cse | and_936_cse
      | and_937_cse;
  assign nor_tmp_230 = while_mux_1418_tmp & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign or_699_nl = and_771_cse | and_770_cse | and_789_cse;
  assign or_697_nl = and_1107_cse | and_1110_cse | nor_tmp_230;
  assign mux_tmp_338 = MUX_s_1_2_2(or_699_nl, or_697_nl, while_stage_0_5);
  assign or_tmp_405 = and_1107_cse | and_1110_cse;
  assign or_tmp_406 = nor_tmp_230 | or_tmp_405;
  assign or_tmp_407 = and_771_cse | and_770_cse;
  assign or_tmp_408 = and_789_cse | or_tmp_407;
  assign nand_18_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_3_sva & (~(weight_mem_read_arbxbar_arbiters_next_3_5_sva
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]))) & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      & (~ or_tmp_407));
  assign mux_342_itm = MUX_s_1_2_2(nand_18_nl, or_tmp_408, and_776_cse);
  assign nand_16_nl = ~(while_mux_1420_tmp & (~(while_mux_1418_tmp & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])))
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]) & (~ or_tmp_405));
  assign mux_340_itm = MUX_s_1_2_2(nand_16_nl, or_tmp_406, and_1108_cse);
  assign mux_345_nl = MUX_s_1_2_2(mux_342_itm, mux_340_itm, while_stage_0_5);
  assign mux_343_nl = MUX_s_1_2_2(mux_342_itm, or_tmp_408, weight_mem_read_arbxbar_arbiters_next_3_1_sva);
  assign mux_341_nl = MUX_s_1_2_2(mux_340_itm, or_tmp_406, while_mux_1422_tmp);
  assign mux_344_nl = MUX_s_1_2_2(mux_343_nl, mux_341_nl, while_stage_0_5);
  assign mux_346_nl = MUX_s_1_2_2(mux_345_nl, mux_344_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign mux_339_nl = MUX_s_1_2_2(or_tmp_408, or_tmp_406, while_stage_0_5);
  assign mux_347_itm = MUX_s_1_2_2(mux_346_nl, mux_339_nl, weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp);
  assign or_708_nl = while_mux_1417_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]));
  assign or_707_nl = while_mux_1416_tmp | and_1107_cse;
  assign mux_348_nl = MUX_s_1_2_2(or_708_nl, or_707_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign mux_349_nl = MUX_s_1_2_2(mux_348_nl, or_tmp_405, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign or_706_nl = while_mux_1418_tmp | or_tmp_405;
  assign mux_350_nl = MUX_s_1_2_2(mux_349_nl, or_706_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign or_tmp_414 = and_1108_cse | mux_350_nl;
  assign or_715_nl = weight_mem_read_arbxbar_arbiters_next_3_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]));
  assign or_714_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1
      | and_771_cse;
  assign mux_351_nl = MUX_s_1_2_2(or_715_nl, or_714_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign mux_352_nl = MUX_s_1_2_2(mux_351_nl, or_tmp_407, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign or_713_nl = weight_mem_read_arbxbar_arbiters_next_3_5_sva | or_tmp_407;
  assign mux_353_nl = MUX_s_1_2_2(mux_352_nl, or_713_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign or_tmp_421 = and_776_cse | mux_353_nl;
  assign mux_358_nl = MUX_s_1_2_2(or_tmp_421, or_tmp_414, while_stage_0_5);
  assign or_721_nl = weight_mem_read_arbxbar_arbiters_next_3_3_sva | or_tmp_421;
  assign or_720_nl = while_mux_1420_tmp | or_tmp_414;
  assign mux_357_nl = MUX_s_1_2_2(or_721_nl, or_720_nl, while_stage_0_5);
  assign mux_359_nl = MUX_s_1_2_2(mux_358_nl, mux_357_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign or_719_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva | or_tmp_421;
  assign or_718_nl = while_mux_1422_tmp | or_tmp_414;
  assign mux_355_nl = MUX_s_1_2_2(or_719_nl, or_718_nl, while_stage_0_5);
  assign or_717_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva | weight_mem_read_arbxbar_arbiters_next_3_3_sva
      | or_tmp_421;
  assign or_710_nl = while_mux_1420_tmp | while_mux_1422_tmp | or_tmp_414;
  assign mux_354_nl = MUX_s_1_2_2(or_717_nl, or_710_nl, while_stage_0_5);
  assign mux_356_nl = MUX_s_1_2_2(mux_355_nl, mux_354_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, mux_356_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign and_dcpl_707 = ~(mux_360_nl | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp);
  assign nor_581_nl = ~(and_776_cse | and_773_cse | and_1106_cse);
  assign nor_582_nl = ~(and_1108_cse | and_1109_cse | and_1111_cse);
  assign mux_361_nl = MUX_s_1_2_2(nor_581_nl, nor_582_nl, while_stage_0_5);
  assign and_dcpl_712 = mux_361_nl & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3])))
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])));
  assign and_1009_cse = while_mux_1410_tmp & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign and_1008_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]) & while_mux_1409_tmp;
  assign or_tmp_442 = and_1008_cse | and_1009_cse;
  assign or_740_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva | or_tmp_442;
  assign or_739_nl = Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 | or_tmp_442;
  assign mux_363_nl = MUX_s_1_2_2(or_740_nl, or_739_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_738_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2])
      | weight_mem_read_arbxbar_arbiters_next_2_5_sva | or_tmp_442;
  assign mux_364_nl = MUX_s_1_2_2(mux_363_nl, or_738_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_365_cse = MUX_s_1_2_2(or_tmp_442, mux_364_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign or_742_nl = and_1114_cse | and_740_cse | and_768_cse;
  assign mux_tmp_366 = MUX_s_1_2_2(or_742_nl, mux_365_cse, while_stage_0_5);
  assign nand_19_nl = ~(while_mux_1412_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      & (~ or_tmp_442));
  assign mux_tmp_370 = MUX_s_1_2_2(nand_19_nl, or_tmp_442, and_1118_cse);
  assign or_752_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva | mux_tmp_370;
  assign or_751_nl = Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 | mux_tmp_370;
  assign mux_371_nl = MUX_s_1_2_2(or_752_nl, or_751_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_750_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2])
      | weight_mem_read_arbxbar_arbiters_next_2_5_sva | mux_tmp_370;
  assign mux_372_nl = MUX_s_1_2_2(mux_371_nl, or_750_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_373 = MUX_s_1_2_2(mux_tmp_370, mux_372_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign or_tmp_459 = and_768_cse | and_740_cse;
  assign or_tmp_460 = and_1114_cse | or_tmp_459;
  assign nand_20_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      & (~ or_tmp_459));
  assign mux_375_nl = MUX_s_1_2_2(nand_20_nl, or_tmp_459, and_767_cse);
  assign or_tmp_461 = and_1114_cse | mux_375_nl;
  assign mux_385_nl = MUX_s_1_2_2(or_tmp_461, mux_tmp_373, while_stage_0_5);
  assign mux_383_nl = MUX_s_1_2_2(or_tmp_461, or_tmp_460, weight_mem_read_arbxbar_arbiters_next_2_2_sva);
  assign mux_382_nl = MUX_s_1_2_2(mux_tmp_373, mux_365_cse, while_mux_1414_tmp);
  assign mux_384_nl = MUX_s_1_2_2(mux_383_nl, mux_382_nl, while_stage_0_5);
  assign mux_386_nl = MUX_s_1_2_2(mux_385_nl, mux_384_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign mux_379_nl = MUX_s_1_2_2(or_tmp_461, or_tmp_460, weight_mem_read_arbxbar_arbiters_next_2_1_sva);
  assign mux_378_nl = MUX_s_1_2_2(mux_tmp_373, mux_365_cse, while_mux_1415_tmp);
  assign mux_380_nl = MUX_s_1_2_2(mux_379_nl, mux_378_nl, while_stage_0_5);
  assign or_753_nl = weight_mem_read_arbxbar_arbiters_next_2_1_sva | weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  assign mux_376_nl = MUX_s_1_2_2(or_tmp_461, or_tmp_460, or_753_nl);
  assign or_743_nl = while_mux_1414_tmp | while_mux_1415_tmp;
  assign mux_374_nl = MUX_s_1_2_2(mux_tmp_373, mux_365_cse, or_743_nl);
  assign mux_377_nl = MUX_s_1_2_2(mux_376_nl, mux_374_nl, while_stage_0_5);
  assign mux_381_nl = MUX_s_1_2_2(mux_380_nl, mux_377_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign mux_387_itm = MUX_s_1_2_2(mux_386_nl, mux_381_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign and_1024_cse = while_mux_1412_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign or_tmp_464 = and_1024_cse | and_1008_cse | and_1009_cse;
  assign and_1034_cse = while_mux_1415_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign and_1028_cse = weight_mem_read_arbxbar_arbiters_next_2_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign mux_393_nl = MUX_s_1_2_2((~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])),
      weight_mem_read_arbxbar_arbiters_next_2_6_sva, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign or_771_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1
      | and_768_cse;
  assign mux_394_nl = MUX_s_1_2_2(mux_393_nl, or_771_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign or_772_nl = and_766_cse | mux_394_nl;
  assign or_770_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva | and_766_cse
      | and_740_cse | and_768_cse;
  assign mux_395_nl = MUX_s_1_2_2(or_772_nl, or_770_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign nor_586_nl = ~(and_767_cse | and_1028_cse | and_738_cse | mux_395_nl);
  assign mux_390_nl = MUX_s_1_2_2((~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])),
      while_mux_1410_tmp, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign or_763_nl = while_mux_1409_tmp | and_1009_cse;
  assign mux_391_nl = MUX_s_1_2_2(mux_390_nl, or_763_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign or_764_nl = and_1024_cse | mux_391_nl;
  assign or_762_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva | or_tmp_464;
  assign or_761_nl = Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 | or_tmp_464;
  assign mux_388_nl = MUX_s_1_2_2(or_762_nl, or_761_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_760_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2])
      | weight_mem_read_arbxbar_arbiters_next_2_5_sva | or_tmp_464;
  assign mux_389_nl = MUX_s_1_2_2(mux_388_nl, or_760_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_392_nl = MUX_s_1_2_2(or_764_nl, mux_389_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign nor_587_nl = ~(and_1118_cse | and_1034_cse | and_1119_cse | mux_392_nl);
  assign not_tmp_443 = MUX_s_1_2_2(nor_586_nl, nor_587_nl, while_stage_0_5);
  assign or_tmp_481 = and_1024_cse | and_1034_cse;
  assign or_tmp_487 = and_766_cse | and_1028_cse;
  assign nor_588_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_1_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])));
  assign nor_589_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_4_sva | and_1028_cse);
  assign mux_400_nl = MUX_s_1_2_2(nor_588_nl, nor_589_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign nor_590_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_2_sva | or_tmp_487);
  assign mux_401_nl = MUX_s_1_2_2(mux_400_nl, nor_590_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign nor_591_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_3_sva | and_738_cse
      | or_tmp_487);
  assign mux_402_nl = MUX_s_1_2_2(mux_401_nl, nor_591_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign nor_592_nl = ~(while_mux_1415_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])));
  assign nor_593_nl = ~(while_mux_1412_tmp | and_1034_cse);
  assign mux_397_nl = MUX_s_1_2_2(nor_592_nl, nor_593_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign nor_594_nl = ~(while_mux_1414_tmp | or_tmp_481);
  assign mux_398_nl = MUX_s_1_2_2(mux_397_nl, nor_594_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign nor_595_nl = ~(while_mux_1413_tmp | and_1119_cse | or_tmp_481);
  assign mux_399_nl = MUX_s_1_2_2(mux_398_nl, nor_595_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign mux_403_nl = MUX_s_1_2_2(mux_402_nl, mux_399_nl, while_stage_0_5);
  assign and_dcpl_717 = mux_403_nl & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])));
  assign or_tmp_496 = and_1024_cse | and_1008_cse | and_1009_cse | and_1034_cse;
  assign or_tmp_509 = and_795_cse | nor_tmp_29;
  assign nor_tmp_317 = Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign and_1049_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) & Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1;
  assign or_tmp_511 = and_1049_cse | nor_tmp_317;
  assign or_tmp_513 = and_795_cse | nor_tmp_317;
  assign or_811_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | nor_tmp_29;
  assign mux_412_nl = MUX_s_1_2_2(or_tmp_513, or_tmp_511, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign mux_411_nl = MUX_s_1_2_2(or_tmp_509, or_811_cse, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign mux_413_nl = MUX_s_1_2_2(mux_412_nl, mux_411_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_414_nl = MUX_s_1_2_2(or_tmp_509, mux_413_nl, while_stage_0_5);
  assign or_810_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_509;
  assign or_809_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_513;
  assign or_807_nl = Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 | or_tmp_511;
  assign mux_408_nl = MUX_s_1_2_2(or_809_nl, or_807_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_805_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1])
      | weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_509;
  assign mux_409_nl = MUX_s_1_2_2(mux_408_nl, or_805_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_410_nl = MUX_s_1_2_2(or_810_nl, mux_409_nl, while_stage_0_5);
  assign mux_tmp_415 = MUX_s_1_2_2(mux_414_nl, mux_410_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign and_752_cse = weight_mem_read_arbxbar_arbiters_next_1_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign and_764_cse = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign and_759_cse = Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign and_758_cse = Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign nand_24_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      & (~ or_tmp_509));
  assign mux_429_nl = MUX_s_1_2_2(nand_24_nl, or_tmp_509, and_794_cse);
  assign mux_430_nl = MUX_s_1_2_2(mux_429_nl, or_tmp_509, and_793_cse);
  assign mux_431_nl = MUX_s_1_2_2(mux_430_nl, or_tmp_509, and_752_cse);
  assign nor_385_nl = ~(and_792_cse | mux_431_nl);
  assign nand_23_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      & (~ or_tmp_513));
  assign mux_424_nl = MUX_s_1_2_2(nand_23_nl, or_tmp_513, and_794_cse);
  assign mux_425_nl = MUX_s_1_2_2(mux_424_nl, or_tmp_513, and_793_cse);
  assign mux_426_nl = MUX_s_1_2_2(mux_425_nl, or_tmp_513, and_752_cse);
  assign nor_386_nl = ~(and_792_cse | mux_426_nl);
  assign nand_22_nl = ~(Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      & (~ or_tmp_511));
  assign mux_421_nl = MUX_s_1_2_2(nand_22_nl, or_tmp_511, and_758_cse);
  assign mux_422_nl = MUX_s_1_2_2(mux_421_nl, or_tmp_511, and_759_cse);
  assign and_760_nl = Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign mux_423_nl = MUX_s_1_2_2(mux_422_nl, or_tmp_511, and_760_nl);
  assign nor_387_nl = ~((Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]))
      | mux_423_nl);
  assign mux_427_nl = MUX_s_1_2_2(nor_386_nl, nor_387_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nand_21_nl = ~(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) & (~ or_tmp_509));
  assign mux_417_nl = MUX_s_1_2_2(nand_21_nl, or_tmp_509, and_794_cse);
  assign mux_418_nl = MUX_s_1_2_2(mux_417_nl, or_tmp_509, and_793_cse);
  assign mux_419_nl = MUX_s_1_2_2(mux_418_nl, or_tmp_509, and_764_cse);
  assign nor_388_nl = ~(and_792_cse | mux_419_nl);
  assign or_815_nl = (~ Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0)
      | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])
      | nor_tmp_29;
  assign or_812_nl = and_764_cse | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign mux_416_nl = MUX_s_1_2_2(or_815_nl, or_811_cse, or_812_nl);
  assign nor_389_nl = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | mux_416_nl);
  assign mux_420_nl = MUX_s_1_2_2(nor_388_nl, nor_389_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign mux_428_nl = MUX_s_1_2_2(mux_427_nl, mux_420_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign not_tmp_449 = MUX_s_1_2_2(nor_385_nl, mux_428_nl, while_stage_0_5);
  assign nor_tmp_350 = while_mux_1408_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign or_tmp_530 = ((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) & while_mux_1405_tmp)
      | nor_tmp_350;
  assign or_tmp_531 = nor_tmp_29 | or_tmp_530;
  assign or_tmp_532 = and_793_cse | or_tmp_531;
  assign or_tmp_534 = and_794_cse | and_795_cse | or_tmp_532;
  assign or_tmp_536 = nor_tmp_317 | or_tmp_530;
  assign or_tmp_537 = and_759_cse | or_tmp_536;
  assign or_tmp_539 = and_758_cse | and_1049_cse | or_tmp_537;
  assign or_tmp_541 = and_793_cse | or_tmp_536;
  assign or_tmp_543 = and_794_cse | and_795_cse | or_tmp_541;
  assign or_tmp_545 = ((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_4_sva)
      | and_752_cse;
  assign or_tmp_547 = and_793_cse | nor_tmp_29 | or_tmp_545;
  assign or_tmp_549 = and_794_cse | and_795_cse | or_tmp_547;
  assign or_845_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_549;
  assign or_839_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_543;
  assign or_835_nl = Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 | or_tmp_539;
  assign mux_433_nl = MUX_s_1_2_2(or_839_nl, or_835_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_830_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1])
      | weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_534;
  assign mux_434_nl = MUX_s_1_2_2(mux_433_nl, or_830_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_435 = MUX_s_1_2_2(or_845_nl, mux_434_nl, while_stage_0_5);
  assign mux_437_nl = MUX_s_1_2_2(or_tmp_543, or_tmp_539, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_847_nl = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]) | or_tmp_531;
  assign mux_436_nl = MUX_s_1_2_2(or_tmp_534, or_847_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign mux_438_nl = MUX_s_1_2_2(mux_437_nl, mux_436_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_439_nl = MUX_s_1_2_2(or_tmp_549, mux_438_nl, while_stage_0_5);
  assign mux_tmp_440 = MUX_s_1_2_2(mux_439_nl, mux_tmp_435, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign or_877_nl = and_793_cse | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      | (~ (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])) | or_tmp_545;
  assign or_854_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva | or_tmp_547;
  assign mux_447_nl = MUX_s_1_2_2(or_877_nl, or_854_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign or_855_nl = and_794_cse | mux_447_nl;
  assign or_878_nl = and_793_cse | Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 | (~
      (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])) | or_tmp_530;
  assign or_852_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva | or_tmp_541;
  assign mux_444_nl = MUX_s_1_2_2(or_878_nl, or_852_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign or_853_nl = and_794_cse | mux_444_nl;
  assign or_879_nl = and_759_cse | Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 | (~
      (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])) | or_tmp_530;
  assign or_850_nl = Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 | or_tmp_537;
  assign mux_443_nl = MUX_s_1_2_2(or_879_nl, or_850_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign or_851_nl = and_758_cse | mux_443_nl;
  assign mux_445_nl = MUX_s_1_2_2(or_853_nl, or_851_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_880_nl = and_793_cse | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      | (~ (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])) | or_tmp_530;
  assign or_848_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva | or_tmp_532;
  assign mux_441_nl = MUX_s_1_2_2(or_880_nl, or_848_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign or_849_nl = and_794_cse | mux_441_nl;
  assign or_881_nl = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]) | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      | (~ (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])) | or_tmp_530;
  assign mux_442_nl = MUX_s_1_2_2(or_849_nl, or_881_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign mux_446_nl = MUX_s_1_2_2(mux_445_nl, mux_442_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_448_nl = MUX_s_1_2_2(or_855_nl, mux_446_nl, while_stage_0_5);
  assign mux_449_nl = MUX_s_1_2_2(mux_448_nl, mux_tmp_435, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign mux_450_itm = MUX_s_1_2_2(mux_449_nl, mux_tmp_440, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign or_858_nl = while_mux_1408_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]));
  assign or_857_nl = while_mux_1405_tmp | nor_tmp_350;
  assign mux_tmp_451 = MUX_s_1_2_2(or_858_nl, or_857_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign or_862_nl = weight_mem_read_arbxbar_arbiters_next_1_3_sva | or_tmp_530;
  assign mux_452_nl = MUX_s_1_2_2(mux_tmp_451, or_862_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign or_861_nl = weight_mem_read_arbxbar_arbiters_next_1_2_sva | and_793_cse
      | or_tmp_530;
  assign mux_tmp_453 = MUX_s_1_2_2(mux_452_nl, or_861_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign or_870_nl = weight_mem_read_arbxbar_arbiters_next_1_1_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]));
  assign or_869_nl = weight_mem_read_arbxbar_arbiters_next_1_4_sva | and_752_cse;
  assign mux_459_nl = MUX_s_1_2_2(or_870_nl, or_869_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign or_868_nl = weight_mem_read_arbxbar_arbiters_next_1_3_sva | or_tmp_545;
  assign mux_460_nl = MUX_s_1_2_2(mux_459_nl, or_868_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign or_867_nl = weight_mem_read_arbxbar_arbiters_next_1_2_sva | and_793_cse
      | or_tmp_545;
  assign mux_461_nl = MUX_s_1_2_2(mux_460_nl, or_867_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign or_865_nl = Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 | or_tmp_530;
  assign mux_455_nl = MUX_s_1_2_2(mux_tmp_451, or_865_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign or_864_nl = Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 | and_759_cse | or_tmp_530;
  assign mux_456_nl = MUX_s_1_2_2(mux_455_nl, or_864_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign mux_457_nl = MUX_s_1_2_2(mux_tmp_453, mux_456_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_859_nl = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | mux_tmp_451;
  assign mux_454_nl = MUX_s_1_2_2(mux_tmp_453, or_859_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign mux_458_nl = MUX_s_1_2_2(mux_457_nl, mux_454_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_462_nl = MUX_s_1_2_2(mux_461_nl, mux_458_nl, while_stage_0_5);
  assign and_dcpl_720 = (~ mux_462_nl) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]))) & nor_428_cse;
  assign and_dcpl_722 = weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp);
  assign and_dcpl_723 = weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_dcpl_724 = ~(weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign or_dcpl_295 = ~(Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs);
  assign PECore_PushAxiRsp_mux_23_itm_1_mx0c1 = and_dcpl_41 & (~ rva_in_reg_rw_sva_5);
  assign and_576_nl = fsm_output & (~ weight_mem_run_3_for_land_4_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000,
      weight_port_read_out_data_3_15_sva_dfm_1, and_576_nl);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[127:120];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_c = {rva_out_reg_data_119_112_sva_dfm_4_1_7
      , rva_out_reg_data_119_112_sva_dfm_4_1_6_0};
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[119:112];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_a = weight_port_read_out_data_7_1_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[15:8];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_c = weight_port_read_out_data_7_0_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[7:0];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_2_a = weight_port_read_out_data_7_3_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[31:24];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_2_c = weight_port_read_out_data_7_2_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[23:16];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_3_a = weight_port_read_out_data_7_5_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[47:40];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_3_c = weight_port_read_out_data_7_4_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[39:32];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_4_a = weight_port_read_out_data_7_7_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[63:56];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_4_c = weight_port_read_out_data_7_6_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[55:48];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_5_a = weight_port_read_out_data_7_9_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[79:72];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_5_c = weight_port_read_out_data_7_8_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[71:64];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_6_a = weight_port_read_out_data_7_11_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[95:88];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_6_c = weight_port_read_out_data_7_10_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[87:80];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_7_a = weight_port_read_out_data_7_13_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[111:104];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_7_c = weight_port_read_out_data_7_12_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[103:96];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_8_a = weight_port_read_out_data_7_15_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[127:120];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_8_c = weight_port_read_out_data_7_14_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[119:112];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_9_a = MUX_v_8_2_2(({weight_port_read_out_data_0_1_sva_mx0_7
      , weight_port_read_out_data_0_1_sva_mx0_6_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_9_c = {weight_port_read_out_data_0_0_sva_dfm_3_7
      , weight_port_read_out_data_0_0_sva_dfm_3_6_0};
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_10_a = MUX_v_8_2_2(({weight_port_read_out_data_0_3_sva_mx0_7_4
      , weight_port_read_out_data_0_3_sva_mx0_3_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_10_c = MUX_v_8_2_2(({weight_port_read_out_data_0_2_sva_mx0_7
      , weight_port_read_out_data_0_2_sva_mx0_6 , weight_port_read_out_data_0_2_sva_mx0_5_4
      , weight_port_read_out_data_0_2_sva_mx0_3_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_11_a = MUX_v_8_2_2(({weight_port_read_out_data_0_5_sva_mx0_7
      , weight_port_read_out_data_0_5_sva_mx0_6_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_11_c = MUX_v_8_2_2(({weight_port_read_out_data_0_4_sva_mx0_7
      , weight_port_read_out_data_0_4_sva_mx0_6_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_12_a = MUX_v_8_2_2(weight_port_read_out_data_0_7_sva_mx0,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_12_c = MUX_v_8_2_2(weight_port_read_out_data_0_6_sva_dfm_2,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_13_a = MUX_v_8_2_2(weight_port_read_out_data_0_9_sva_dfm_2,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_13_c = MUX_v_8_2_2(weight_port_read_out_data_0_8_sva_dfm_2,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_14_a = MUX_v_8_2_2(({weight_port_read_out_data_0_11_sva_dfm_2_7
      , weight_port_read_out_data_0_11_sva_dfm_2_6 , weight_port_read_out_data_0_11_sva_dfm_2_5_4
      , weight_port_read_out_data_0_11_sva_dfm_2_3_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_14_c = MUX_v_8_2_2(({weight_port_read_out_data_0_10_sva_dfm_2_7
      , weight_port_read_out_data_0_10_sva_dfm_2_6_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_15_a = MUX_v_8_2_2(({weight_port_read_out_data_0_13_sva_dfm_2_7
      , weight_port_read_out_data_0_13_sva_dfm_2_6_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_15_c = MUX_v_8_2_2(({weight_port_read_out_data_0_12_sva_dfm_2_7_4
      , weight_port_read_out_data_0_12_sva_dfm_2_3_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_16_a = MUX_v_8_2_2(weight_port_read_out_data_0_15_sva_dfm_2,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_16_c = MUX_v_8_2_2(({weight_port_read_out_data_0_14_sva_dfm_2_7
      , weight_port_read_out_data_0_14_sva_dfm_2_6_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_17_a = MUX_v_8_2_2(weight_port_read_out_data_6_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_17_c = MUX_v_8_2_2(weight_port_read_out_data_6_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_18_a = MUX_v_8_2_2(weight_port_read_out_data_6_3_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_18_c = MUX_v_8_2_2(weight_port_read_out_data_6_2_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_19_a = MUX_v_8_2_2(weight_port_read_out_data_6_5_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_19_c = MUX_v_8_2_2(weight_port_read_out_data_6_4_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_20_a = MUX_v_8_2_2(weight_port_read_out_data_6_7_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_20_c = MUX_v_8_2_2(weight_port_read_out_data_6_6_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_21_a = MUX_v_8_2_2(weight_port_read_out_data_6_9_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_21_c = MUX_v_8_2_2(weight_port_read_out_data_6_8_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_22_a = MUX_v_8_2_2(weight_port_read_out_data_6_11_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_22_c = MUX_v_8_2_2(weight_port_read_out_data_6_10_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_23_a = MUX_v_8_2_2(weight_port_read_out_data_6_13_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_23_c = MUX_v_8_2_2(weight_port_read_out_data_6_12_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_24_a = MUX_v_8_2_2(weight_port_read_out_data_6_15_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_24_c = MUX_v_8_2_2(weight_port_read_out_data_6_14_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_25_a = MUX_v_8_2_2(weight_port_read_out_data_1_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_25_c = MUX_v_8_2_2(weight_port_read_out_data_1_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_26_a = MUX_v_8_2_2(weight_port_read_out_data_1_3_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_26_c = MUX_v_8_2_2(weight_port_read_out_data_1_2_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_27_a = MUX_v_8_2_2(weight_port_read_out_data_1_5_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_27_c = MUX_v_8_2_2(weight_port_read_out_data_1_4_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_28_a = MUX_v_8_2_2(weight_port_read_out_data_1_7_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_28_c = MUX_v_8_2_2(weight_port_read_out_data_1_6_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_29_a = MUX_v_8_2_2(weight_port_read_out_data_1_9_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_29_c = MUX_v_8_2_2(weight_port_read_out_data_1_8_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_30_a = MUX_v_8_2_2(weight_port_read_out_data_1_11_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_30_c = MUX_v_8_2_2(weight_port_read_out_data_1_10_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_31_a = MUX_v_8_2_2(weight_port_read_out_data_1_13_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_31_c = MUX_v_8_2_2(weight_port_read_out_data_1_12_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign and_575_nl = fsm_output & (~ weight_mem_run_3_for_land_2_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_32_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000,
      weight_port_read_out_data_1_15_sva_dfm_1, and_575_nl);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_32_c = {rva_out_reg_data_103_96_sva_dfm_4_1_7_4
      , rva_out_reg_data_103_96_sva_dfm_4_1_3_0};
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_33_a = MUX_v_8_2_2(weight_port_read_out_data_5_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_33_c = MUX_v_8_2_2(weight_port_read_out_data_5_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_34_a = MUX_v_8_2_2(weight_port_read_out_data_5_3_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_34_c = MUX_v_8_2_2(weight_port_read_out_data_5_2_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_35_a = MUX_v_8_2_2(weight_port_read_out_data_5_5_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_35_c = MUX_v_8_2_2(weight_port_read_out_data_5_4_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_36_a = MUX_v_8_2_2(weight_port_read_out_data_5_7_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_36_c = MUX_v_8_2_2(weight_port_read_out_data_5_6_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_37_a = MUX_v_8_2_2(weight_port_read_out_data_5_9_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_37_c = MUX_v_8_2_2(weight_port_read_out_data_5_8_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_38_a = MUX_v_8_2_2(weight_port_read_out_data_5_11_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_38_c = MUX_v_8_2_2(weight_port_read_out_data_5_10_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_39_a = MUX_v_8_2_2(weight_port_read_out_data_5_13_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_39_c = MUX_v_8_2_2(weight_port_read_out_data_5_12_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
      weight_mem_run_3_for_land_6_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_40_a = weight_port_read_out_data_5_15_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_40_c = weight_port_read_out_data_5_14_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_41_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_port_read_out_data_2_1_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_41_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[15:8];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_41_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
      weight_port_read_out_data_2_0_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_41_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[7:0];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_42_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
      weight_port_read_out_data_2_3_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_42_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[31:24];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_42_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
      weight_port_read_out_data_2_2_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_42_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[23:16];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_43_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
      weight_port_read_out_data_2_5_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_43_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[47:40];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_43_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
      weight_port_read_out_data_2_4_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_43_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[39:32];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_44_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
      weight_port_read_out_data_2_7_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_44_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[63:56];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_44_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
      weight_port_read_out_data_2_6_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_44_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[55:48];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_45_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
      weight_port_read_out_data_2_9_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_45_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[79:72];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_45_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
      weight_port_read_out_data_2_8_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_45_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[71:64];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_46_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
      weight_port_read_out_data_2_11_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_46_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[95:88];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_46_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
      weight_port_read_out_data_2_10_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_46_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[87:80];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_47_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
      weight_port_read_out_data_2_13_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_47_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[111:104];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_47_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
      weight_port_read_out_data_2_12_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_47_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[103:96];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_48_a = {rva_out_reg_data_111_104_sva_dfm_4_1_7
      , rva_out_reg_data_111_104_sva_dfm_4_1_6_0};
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_48_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014,
      weight_port_read_out_data_2_14_sva_dfm_1, and_dcpl_562);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_49_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_port_read_out_data_4_1_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_49_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
      weight_port_read_out_data_4_0_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_50_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
      weight_port_read_out_data_4_3_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_50_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
      weight_port_read_out_data_4_2_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_51_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
      weight_port_read_out_data_4_5_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_51_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
      weight_port_read_out_data_4_4_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_52_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
      weight_port_read_out_data_4_7_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_52_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
      weight_port_read_out_data_4_6_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_53_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
      weight_port_read_out_data_4_9_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_53_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
      weight_port_read_out_data_4_8_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_54_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
      weight_port_read_out_data_4_11_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_54_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
      weight_port_read_out_data_4_10_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_55_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
      weight_port_read_out_data_4_13_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_55_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
      weight_port_read_out_data_4_12_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_56_a = rva_out_reg_data_127_120_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_56_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014,
      weight_port_read_out_data_4_14_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_57_a = MUX_v_8_2_2(weight_port_read_out_data_3_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_57_c = MUX_v_8_2_2(weight_port_read_out_data_3_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_58_a = MUX_v_8_2_2(weight_port_read_out_data_3_3_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_58_c = MUX_v_8_2_2(weight_port_read_out_data_3_2_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_59_a = MUX_v_8_2_2(weight_port_read_out_data_3_5_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_59_c = MUX_v_8_2_2(weight_port_read_out_data_3_4_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_60_a = MUX_v_8_2_2(weight_port_read_out_data_3_7_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_60_c = MUX_v_8_2_2(weight_port_read_out_data_3_6_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_61_a = MUX_v_8_2_2(weight_port_read_out_data_3_9_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_61_c = MUX_v_8_2_2(weight_port_read_out_data_3_8_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_62_a = MUX_v_8_2_2(weight_port_read_out_data_3_11_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_62_c = MUX_v_8_2_2(weight_port_read_out_data_3_10_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_63_a = MUX_v_8_2_2(weight_port_read_out_data_3_13_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_63_c = MUX_v_8_2_2(weight_port_read_out_data_3_12_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0));
  assign weight_mem_banks_write_if_for_if_and_35_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_36_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_37_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_38_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_39_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_40_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_41_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      , weight_mem_banks_write_if_for_if_and_35_nl , weight_mem_banks_write_if_for_if_and_36_nl
      , weight_mem_banks_write_if_for_if_and_37_nl , weight_mem_banks_write_if_for_if_and_38_nl
      , weight_mem_banks_write_if_for_if_and_39_nl , weight_mem_banks_write_if_for_if_and_40_nl
      , weight_mem_banks_write_if_for_if_and_41_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0});
  assign weight_mem_banks_write_if_for_if_mux_7_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      , weight_mem_banks_write_if_for_if_mux_7_nl};
  assign nor_610_nl = ~((~ PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3) |
      PECore_RunFSM_switch_lp_equal_tmp_1_2);
  assign mux_159_nl = MUX_s_1_2_2(or_79_cse, nor_610_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff = mux_159_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_2[14:3];
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff = and_dcpl_189;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0));
  assign weight_mem_banks_write_if_for_if_and_28_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_29_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_30_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_31_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_32_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_33_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_34_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      , weight_mem_banks_write_if_for_if_and_28_nl , weight_mem_banks_write_if_for_if_and_29_nl
      , weight_mem_banks_write_if_for_if_and_30_nl , weight_mem_banks_write_if_for_if_and_31_nl
      , weight_mem_banks_write_if_for_if_and_32_nl , weight_mem_banks_write_if_for_if_and_33_nl
      , weight_mem_banks_write_if_for_if_and_34_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0});
  assign weight_mem_banks_write_if_for_if_mux_6_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      , weight_mem_banks_write_if_for_if_mux_6_nl};
  assign nor_609_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ mux_tmp_130));
  assign mux_158_nl = MUX_s_1_2_2(mux_tmp_131, nor_609_nl, PECore_UpdateFSM_switch_lp_equal_tmp_2_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff = mux_158_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff = and_dcpl_192;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0));
  assign weight_mem_banks_write_if_for_if_and_21_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_22_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_23_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_24_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_25_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_26_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_27_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      , weight_mem_banks_write_if_for_if_and_21_nl , weight_mem_banks_write_if_for_if_and_22_nl
      , weight_mem_banks_write_if_for_if_and_23_nl , weight_mem_banks_write_if_for_if_and_24_nl
      , weight_mem_banks_write_if_for_if_and_25_nl , weight_mem_banks_write_if_for_if_and_26_nl
      , weight_mem_banks_write_if_for_if_and_27_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0});
  assign weight_mem_banks_write_if_for_if_mux_5_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      , weight_mem_banks_write_if_for_if_mux_5_nl};
  assign nor_608_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_3) | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]));
  assign mux_157_nl = MUX_s_1_2_2(mux_tmp_126, nor_608_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff = mux_157_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff = and_dcpl_195;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0));
  assign weight_mem_banks_write_if_for_if_and_14_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_15_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_16_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_17_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_18_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_19_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_20_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      , weight_mem_banks_write_if_for_if_and_14_nl , weight_mem_banks_write_if_for_if_and_15_nl
      , weight_mem_banks_write_if_for_if_and_16_nl , weight_mem_banks_write_if_for_if_and_17_nl
      , weight_mem_banks_write_if_for_if_and_18_nl , weight_mem_banks_write_if_for_if_and_19_nl
      , weight_mem_banks_write_if_for_if_and_20_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0});
  assign weight_mem_banks_write_if_for_if_mux_4_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      , weight_mem_banks_write_if_for_if_mux_4_nl};
  assign nor_607_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3) | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]));
  assign mux_156_nl = MUX_s_1_2_2(or_100_cse, nor_607_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff = mux_156_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff = and_dcpl_545;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0));
  assign weight_mem_banks_write_if_for_if_and_7_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_9_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_10_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_11_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_12_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_13_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      , weight_mem_banks_write_if_for_if_and_7_nl , weight_mem_banks_write_if_for_if_and_8_nl
      , weight_mem_banks_write_if_for_if_and_9_nl , weight_mem_banks_write_if_for_if_and_10_nl
      , weight_mem_banks_write_if_for_if_and_11_nl , weight_mem_banks_write_if_for_if_and_12_nl
      , weight_mem_banks_write_if_for_if_and_13_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0});
  assign weight_mem_banks_write_if_for_if_mux_3_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      , weight_mem_banks_write_if_for_if_mux_3_nl};
  assign nor_606_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1)
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]));
  assign mux_155_nl = MUX_s_1_2_2(or_tmp_136, nor_606_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff = mux_155_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff = and_dcpl_200;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0));
  assign weight_mem_banks_write_if_for_if_and_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_1_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_2_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_3_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_5_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl ,
      weight_mem_banks_write_if_for_if_and_nl , weight_mem_banks_write_if_for_if_and_1_nl
      , weight_mem_banks_write_if_for_if_and_2_nl , weight_mem_banks_write_if_for_if_and_3_nl
      , weight_mem_banks_write_if_for_if_and_4_nl , weight_mem_banks_write_if_for_if_and_5_nl
      , weight_mem_banks_write_if_for_if_and_6_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0});
  assign weight_mem_banks_write_if_for_if_mux_2_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      , weight_mem_banks_write_if_for_if_mux_2_nl};
  assign nor_605_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1)
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]));
  assign mux_154_nl = MUX_s_1_2_2(mux_tmp_115, nor_605_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff = mux_154_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff = and_dcpl_202;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_14_lpi_1_dfm_1_3_2 , weight_write_data_data_0_13_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_12_lpi_1_dfm_1_3_2 , weight_write_data_data_0_11_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_10_lpi_1_dfm_1_3_2 , weight_write_data_data_0_9_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_8_lpi_1_dfm_1_3_2 , weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_1_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_54_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0,
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_1_nl
      , weight_mem_banks_write_if_for_if_mux_54_nl};
  assign nor_604_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1);
  assign mux_153_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_604_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff = mux_153_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_3_14_3;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff = and_dcpl_537;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_14_lpi_1_dfm_1_3_2 , weight_write_data_data_0_13_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_12_lpi_1_dfm_1_3_2 , weight_write_data_data_0_11_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_10_lpi_1_dfm_1_3_2 , weight_write_data_data_0_9_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_8_lpi_1_dfm_1_3_2 , weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_53_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0,
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_nl
      , weight_mem_banks_write_if_for_if_mux_53_nl};
  assign nor_603_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1);
  assign mux_152_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_603_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff = mux_152_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff = and_dcpl_534;
  assign and_dcpl = (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1;
  assign and_dcpl_725 = (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1;
  assign or_dcpl = and_dcpl_725 | and_dcpl;
  assign or_dcpl_296 = and_dcpl_725 | ((pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1);
  assign or_dcpl_298 = ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]) & nor_436_cse)
      | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]) & and_dcpl_657) | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1])
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]));
  assign or_dcpl_300 = ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]) & and_dcpl_662)
      | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]) & and_dcpl_661) | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1])
      & and_dcpl_659);
  assign or_dcpl_301 = ((~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1])) &
      (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]) & and_dcpl_663)
      | (and_dcpl_670 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign and_dcpl_737 = or_dcpl_298 & and_dcpl_663;
  assign and_676_ssc = and_dcpl_663 & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign and_677_ssc = and_dcpl_663 & and_dcpl_657;
  assign and_678_ssc = and_dcpl_663 & nor_436_cse;
  assign and_680_ssc = (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      & weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_683_ssc = and_dcpl_670 & (~(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4));
  assign and_686_ssc = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign PECore_DecodeAxiRead_switch_lp_mux_21_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[0]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl
      = PECore_DecodeAxiRead_switch_lp_mux_21_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_36_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl,
      rva_out_reg_data_0_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_24_itm = MUX_s_1_2_2(rva_out_reg_data_mux_36_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_DecodeAxiRead_switch_lp_mux_22_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[8]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl
      = PECore_DecodeAxiRead_switch_lp_mux_22_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_37_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl,
      rva_out_reg_data_8_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_25_itm = MUX_s_1_2_2(rva_out_reg_data_mux_37_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_DecodeAxiRead_switch_lp_mux_23_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[16]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl
      = PECore_DecodeAxiRead_switch_lp_mux_23_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_38_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl,
      rva_out_reg_data_16_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_26_itm = MUX_s_1_2_2(rva_out_reg_data_mux_38_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_DecodeAxiRead_switch_lp_mux_24_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[24]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl
      = PECore_DecodeAxiRead_switch_lp_mux_24_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_40_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl,
      rva_out_reg_data_24_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_27_nl = MUX_s_1_2_2(rva_out_reg_data_mux_40_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_PushAxiRsp_if_mux1h_15 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_27_nl,
      (weight_port_read_out_data_0_3_sva_dfm_5_rsp_1[0]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl
      = (SC_SRAM_CONFIG[31]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9) &
      PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_39_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl,
      rva_out_reg_data_31_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_28_nl = MUX_s_1_2_2(rva_out_reg_data_mux_39_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_PushAxiRsp_if_mux1h_17 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_28_nl,
      (weight_port_read_out_data_0_3_sva_dfm_5_rsp_0[3]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign weight_port_read_out_data_and_131_ssc = PECoreRun_wen & (~(mux_6_itm & (~((~
      rva_in_reg_rw_sva_st_1_5) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3))
      & while_stage_0_6)) & and_dcpl_41;
  assign and_1624_cse = weight_mem_run_3_for_land_1_lpi_1_dfm_2 & while_stage_0_6;
  assign and_1625_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & while_stage_0_6;
  assign mux_567_nl = MUX_s_1_2_2((~ mux_565_cse), or_tmp_623, and_1624_cse);
  assign mux_566_nl = MUX_s_1_2_2((~ mux_565_cse), or_tmp_623, and_1625_cse);
  assign mux_568_nl = MUX_s_1_2_2(mux_567_nl, mux_566_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_1562_cse = (~ mux_568_nl) & and_dcpl_41 & PECoreRun_wen;
  assign and_1155_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_dcpl_296);
  assign mux_32_nl = MUX_s_1_2_2(or_tmp_47, mux_tmp_31, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign weight_mem_banks_load_store_for_else_and_56_ssc = PECoreRun_wen & (~ mux_32_nl)
      & and_dcpl_48;
  assign or_211_nl = rva_in_reg_rw_sva_st_4 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 | rva_in_reg_rw_sva_4 | (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3)
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1
      | rva_in_reg_rw_sva_st_1_4;
  assign mux_34_nl = MUX_s_1_2_2(or_211_nl, mux_tmp_31, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign weight_mem_banks_load_store_for_else_and_68_ssc = PECoreRun_wen & (~ mux_34_nl)
      & and_dcpl_48;
  assign nor_494_nl = ~((~((~((~((~((~(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign nor_495_nl = ~(rva_in_reg_rw_sva_st_1_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1
      | rva_in_reg_rw_sva_st_4 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4
      | rva_in_reg_rw_sva_4 | (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3) |
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4);
  assign mux_35_nl = MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]),
      (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign nor_496_nl = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2])
      | (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]));
  assign mux_36_nl = MUX_s_1_2_2(mux_35_nl, nor_496_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_37_nl = MUX_s_1_2_2(nor_495_nl, mux_36_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_38_nl = MUX_s_1_2_2(nor_494_nl, mux_37_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_load_store_for_else_and_75_ssc = PECoreRun_wen & mux_38_nl
      & while_stage_0_6;
  assign weight_port_read_out_data_and_225_enex5 = weight_port_read_out_data_and_182_ssc
      & reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo;
  assign weight_port_read_out_data_and_185_ssc = PECoreRun_wen & and_dcpl_279 & (~
      rva_in_reg_rw_sva_st_1_6) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
  assign weight_port_read_out_data_and_226_enex5 = weight_port_read_out_data_and_185_ssc
      & reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo_1;
  assign weight_port_read_out_data_and_227_enex5 = weight_port_read_out_data_and_185_ssc
      & reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo;
  assign weight_port_read_out_data_and_228_enex5 = weight_port_read_out_data_and_185_ssc
      & reg_weight_port_read_out_data_0_2_sva_dfm_1_2_enexo;
  assign weight_port_read_out_data_and_229_enex5 = weight_port_read_out_data_and_185_ssc
      & reg_weight_port_read_out_data_0_3_sva_dfm_1_enexo;
  assign weight_port_read_out_data_and_230_enex5 = weight_port_read_out_data_and_185_ssc
      & reg_weight_port_read_out_data_0_3_sva_dfm_1_1_enexo;
  assign or_306_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign weight_port_read_out_data_and_189_ssc = PECoreRun_wen & and_dcpl_403 & or_306_cse;
  assign and_1183_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_894_tmp);
  assign and_1184_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_1_cse & (~
      or_894_tmp);
  assign and_1185_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      & (~ or_894_tmp);
  assign and_1186_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1
      & (~ or_894_tmp);
  assign and_1187_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      & (~ or_894_tmp);
  assign and_1188_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      & (~ or_894_tmp);
  assign nor_630_ssc = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_894_tmp);
  assign mux1h_5_nl = MUX1HOT_s_1_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[47]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[47]),
      weight_port_read_out_data_0_5_sva_mx0_7, {and_1183_ssc , and_1184_ssc , and_1185_ssc
      , and_1186_ssc , and_1187_ssc , and_1188_ssc , nor_630_ssc});
  assign weight_port_read_out_data_0_5_sva_dfm_mx0w2_7 = mux1h_5_nl & (~ or_894_tmp);
  assign mux1h_12_nl = MUX1HOT_v_7_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[46:40]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[46:40]),
      weight_port_read_out_data_0_5_sva_mx0_6_0, {and_1183_ssc , and_1184_ssc , and_1185_ssc
      , and_1186_ssc , and_1187_ssc , and_1188_ssc , nor_630_ssc});
  assign not_2450_nl = ~ or_894_tmp;
  assign weight_port_read_out_data_0_5_sva_dfm_mx0w2_6_0 = MUX_v_7_2_2(7'b0000000,
      mux1h_12_nl, not_2450_nl);
  assign and_1191_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 & (~ or_dcpl);
  assign and_1193_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      & (~ or_dcpl);
  assign and_1194_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      & (~ or_dcpl);
  assign mux1h_6_nl = MUX1HOT_s_1_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[39]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[39]),
      weight_port_read_out_data_0_4_sva_mx0_7, {and_1191_ssc , and_1148_cse , and_1193_ssc
      , and_1194_ssc , and_1151_cse , and_1152_cse , nor_626_cse});
  assign weight_port_read_out_data_0_4_sva_dfm_mx0w2_7 = mux1h_6_nl & (~ or_dcpl);
  assign mux1h_13_nl = MUX1HOT_v_7_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[38:32]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[38:32]),
      weight_port_read_out_data_0_4_sva_mx0_6_0, {and_1191_ssc , and_1148_cse , and_1193_ssc
      , and_1194_ssc , and_1151_cse , and_1152_cse , nor_626_cse});
  assign not_2451_nl = ~ or_dcpl;
  assign weight_port_read_out_data_0_4_sva_dfm_mx0w2_6_0 = MUX_v_7_2_2(7'b0000000,
      mux1h_13_nl, not_2451_nl);
  assign and_1199_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 & (~ or_dcpl_296);
  assign mux1h_7_nl = MUX1HOT_s_1_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[7]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[7]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[7]),
      weight_port_read_out_data_0_0_sva_dfm_2_7_1, {and_1199_ssc , and_1156_cse ,
      and_1157_cse , and_1158_cse , and_1159_cse , and_1160_cse , nor_627_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w0_7 = mux1h_7_nl & (~ or_dcpl_296);
  assign mux1h_14_nl = MUX1HOT_v_7_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_6_0,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[6:0]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[6:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[6:0]),
      weight_port_read_out_data_0_0_sva_dfm_2_6_0_1, {and_1199_ssc , and_1156_cse
      , and_1157_cse , and_1158_cse , and_1159_cse , and_1160_cse , nor_627_cse});
  assign not_2452_nl = ~ or_dcpl_296;
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w0_6_0 = MUX_v_7_2_2(7'b0000000,
      mux1h_14_nl, not_2452_nl);
  assign weight_port_read_out_data_and_231_enex5 = weight_port_read_out_data_and_123_cse
      & reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_1_enexo;
  assign weight_port_read_out_data_and_232_enex5 = weight_port_read_out_data_and_123_cse
      & reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_1_enexo;
  assign weight_port_read_out_data_and_233_enex5 = weight_port_read_out_data_and_123_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_4_enexo;
  assign weight_port_read_out_data_and_234_enex5 = weight_port_read_out_data_and_123_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_4_1_enexo;
  assign mux_5_nl = MUX_s_1_2_2(and_1619_cse, mux_tmp_4, while_stage_0_7);
  assign weight_port_read_out_data_and_130_ssc = PECoreRun_wen & mux_5_nl;
  assign nor_743_nl = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_2 | (~ mux_tmp_546));
  assign mux_591_nl = MUX_s_1_2_2(mux_tmp_546, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_592_nl = MUX_s_1_2_2(nor_743_nl, mux_591_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_593_nl = MUX_s_1_2_2(mux_tmp_546, mux_592_nl, while_stage_0_6);
  assign and_1578_cse = mux_593_nl & PECoreRun_wen;
  assign weight_port_read_out_data_and_235_enex5 = weight_port_read_out_data_and_174_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo;
  assign weight_port_read_out_data_and_236_enex5 = weight_port_read_out_data_and_174_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_3_enexo;
  assign weight_port_read_out_data_and_237_enex5 = weight_port_read_out_data_and_174_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_3_1_enexo;
  assign weight_port_read_out_data_0_0_sva_dfm_3_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_0_sva_dfm_2_7_1,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[7]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[7]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_145_cse
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , weight_mem_run_3_for_5_and_148_itm_2 , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , weight_mem_run_3_for_5_and_150_itm_2 , reg_weight_mem_run_3_for_5_and_151_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_3_6_0 = MUX1HOT_v_7_9_2(weight_port_read_out_data_0_0_sva_dfm_2_6_0_1,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[6:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[6:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[6:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[6:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[6:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[6:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[6:0]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[6:0]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_145_cse
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , weight_mem_run_3_for_5_and_148_itm_2 , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , weight_mem_run_3_for_5_and_150_itm_2 , reg_weight_mem_run_3_for_5_and_151_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign weight_port_read_out_data_0_5_sva_mx0_7 = MUX1HOT_s_1_3_2(weight_port_read_out_data_0_2_sva_dfm_1_1_7,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7,
      weight_port_read_out_data_0_5_sva_rsp_0, {and_dcpl_279 , and_dcpl_277 , (~
      while_stage_0_8)});
  assign weight_port_read_out_data_0_5_sva_mx0_6_0 = MUX1HOT_v_7_3_2(({weight_port_read_out_data_0_2_sva_dfm_1_1_6
      , weight_port_read_out_data_0_2_sva_dfm_1_1_5_4 , weight_port_read_out_data_0_2_sva_dfm_1_1_3_0}),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0,
      weight_port_read_out_data_0_5_sva_rsp_1, {and_dcpl_279 , and_dcpl_277 , (~
      while_stage_0_8)});
  assign weight_port_read_out_data_0_4_sva_mx0_7 = MUX1HOT_s_1_3_2(weight_port_read_out_data_0_1_sva_dfm_1_1_7,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7,
      weight_port_read_out_data_0_4_sva_rsp_0, {and_dcpl_279 , and_dcpl_277 , (~
      while_stage_0_8)});
  assign weight_port_read_out_data_0_4_sva_mx0_6_0 = MUX1HOT_v_7_3_2(weight_port_read_out_data_0_1_sva_dfm_1_1_6_0,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0,
      weight_port_read_out_data_0_4_sva_rsp_1, {and_dcpl_279 , and_dcpl_277 , (~
      while_stage_0_8)});
  assign weight_port_read_out_data_0_3_sva_mx0_7_4 = MUX1HOT_v_4_3_2(weight_port_read_out_data_0_3_sva_dfm_1_7_4,
      weight_port_read_out_data_0_3_sva_dfm_1_1_7_4, weight_port_read_out_data_0_3_sva_7_4,
      {and_dcpl_279 , and_dcpl_277 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_3_sva_mx0_3_0 = MUX1HOT_v_4_3_2(weight_port_read_out_data_0_3_sva_dfm_1_3_0,
      weight_port_read_out_data_0_3_sva_dfm_1_1_3_0, weight_port_read_out_data_0_3_sva_3_0,
      {and_dcpl_279 , and_dcpl_277 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_2_sva_mx0_7 = MUX1HOT_s_1_3_2(weight_port_read_out_data_0_2_sva_dfm_1_7,
      weight_port_read_out_data_0_2_sva_dfm_1_1_7, reg_weight_port_read_out_data_0_2_ftd,
      {and_dcpl_279 , and_dcpl_277 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_2_sva_mx0_6 = MUX1HOT_s_1_3_2(weight_port_read_out_data_0_2_sva_dfm_1_6,
      weight_port_read_out_data_0_2_sva_dfm_1_1_6, reg_weight_port_read_out_data_0_2_ftd_1,
      {and_dcpl_279 , and_dcpl_277 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_2_sva_mx0_5_4 = MUX1HOT_v_2_3_2(weight_port_read_out_data_0_2_sva_dfm_1_5_4,
      weight_port_read_out_data_0_2_sva_dfm_1_1_5_4, weight_port_read_out_data_0_2_sva_5_4,
      {and_dcpl_279 , and_dcpl_277 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_2_sva_mx0_3_0 = MUX1HOT_v_4_3_2(weight_port_read_out_data_0_2_sva_dfm_1_3_0,
      weight_port_read_out_data_0_2_sva_dfm_1_1_3_0, weight_port_read_out_data_0_2_sva_3_0,
      {and_dcpl_279 , and_dcpl_277 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_1_sva_mx0_7 = MUX1HOT_s_1_3_2(weight_port_read_out_data_0_1_sva_dfm_1_7,
      weight_port_read_out_data_0_1_sva_dfm_1_1_7, weight_port_read_out_data_0_1_sva_7,
      {and_dcpl_279 , and_dcpl_277 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_1_sva_mx0_6_0 = MUX1HOT_v_7_3_2(weight_port_read_out_data_0_1_sva_dfm_1_6_0,
      weight_port_read_out_data_0_1_sva_dfm_1_1_6_0, weight_port_read_out_data_0_1_sva_6_0,
      {and_dcpl_279 , and_dcpl_277 , (~ while_stage_0_8)});
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1_3 = MUX_s_1_2_2(rva_out_reg_data_39_36_sva_dfm_4_1_3,
      rva_out_reg_data_39_36_sva_dfm_6_rsp_0, or_dcpl_291);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1_2_0 = MUX_v_3_2_2(rva_out_reg_data_39_36_sva_dfm_4_1_2_0,
      rva_out_reg_data_39_36_sva_dfm_6_rsp_1, or_dcpl_291);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_107_nl
      = (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[95]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]));
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_123_nl
      = (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[95]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1_7
      = MUX_s_1_8_2(weight_port_read_out_data_0_2_sva_dfm_1_1_7, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_107_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_123_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_106_nl
      = (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[87]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]));
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_122_nl
      = (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[87]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_sva_1_7
      = MUX_s_1_8_2(weight_port_read_out_data_0_1_sva_dfm_1_1_7, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_106_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_122_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_275_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_133_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[86:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_275_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_276_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_134_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[86:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_276_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000000
      = MUX_v_7_8_2(weight_port_read_out_data_0_1_sva_dfm_1_1_6_0, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_133_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_134_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign rva_out_reg_data_and_214_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_1_1_enexo;
  assign while_if_while_if_and_27_nl = MUX_v_4_2_2(4'b0000, rva_out_reg_data_103_96_sva_dfm_6_7_4,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_103_96_sva_dfm_4_mx0w0_7_4 = MUX1HOT_v_4_3_2(while_if_while_if_and_27_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:100]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_s000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_35_nl = MUX_v_4_2_2(4'b0000, rva_out_reg_data_103_96_sva_dfm_6_3_0,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_103_96_sva_dfm_4_mx0w0_3_0 = MUX1HOT_v_4_3_2(while_if_while_if_and_35_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[99:96]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_s000001,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_95_88_sva_dfm_7_7 = MUX1HOT_s_1_3_2(rva_out_reg_data_95_88_sva_dfm_8_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[95]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1_7,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_95_88_sva_dfm_7_6 = MUX1HOT_s_1_3_2(rva_out_reg_data_95_88_sva_dfm_8_6,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[94]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1_6,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_95_88_sva_dfm_7_5_4 = MUX1HOT_v_2_3_2(rva_out_reg_data_95_88_sva_dfm_8_5_4,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[93:92]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_s000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_37_nl = MUX_v_4_2_2(4'b0000, rva_out_reg_data_95_88_sva_dfm_6_3_0,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_95_88_sva_dfm_7_3_0 = MUX1HOT_v_4_3_2(while_if_while_if_and_37_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[91:88]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_s000001,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_87_80_sva_dfm_7_7 = MUX1HOT_s_1_3_2(rva_out_reg_data_87_80_sva_dfm_8_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[87]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_sva_1_7,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_33_nl = MUX_v_7_2_2(7'b0000000, rva_out_reg_data_87_80_sva_dfm_6_6_0,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_87_80_sva_dfm_7_6_0 = MUX1HOT_v_7_3_2(while_if_while_if_and_33_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[86:80]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_110_nl
      = (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[119]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]));
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_126_nl
      = (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[119]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000
      = MUX_s_1_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_110_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_126_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_281_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_145_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[118:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_281_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_282_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_146_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[118:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_282_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001
      = MUX_v_7_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_145_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_146_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_109_nl
      = (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[111]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]));
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_125_nl
      = (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[111]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000
      = MUX_s_1_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_109_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_125_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_283_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_147_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[110:104]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_283_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_284_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_148_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[110:104]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_284_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001
      = MUX_v_7_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_147_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_148_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_279_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_108_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[103:100]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_279_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_280_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_124_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[103:100]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_280_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_s000000
      = MUX_v_4_8_2(weight_port_read_out_data_0_3_sva_dfm_1_1_7_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_108_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_124_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_147_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_139_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[99:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_147_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_162_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_140_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[99:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_162_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_s000001
      = MUX_v_4_8_2(weight_port_read_out_data_0_3_sva_dfm_1_1_3_0, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_139_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_140_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl
      = (SC_SRAM_CONFIG[7]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9) &
      PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_10_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl,
      rva_out_reg_data_7_1_sva_dfm_6_6, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5[6]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_6, {PECore_PushAxiRsp_if_asn_79
      , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl
      = (SC_SRAM_CONFIG[6:1]) & (signext_6_1(~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9))
      & ({{5{PECore_DecodeAxiRead_switch_lp_nor_9_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1});
  assign PECore_PushAxiRsp_if_mux1h_10_5_0 = MUX1HOT_v_6_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl,
      rva_out_reg_data_7_1_sva_dfm_6_5_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5[5:0]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_5_0,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_18_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[15]),
      (rva_out_reg_data_15_9_sva_dfm_10[6]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl
      = PECore_DecodeAxiRead_switch_lp_mux_18_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_12_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl,
      rva_out_reg_data_15_9_sva_dfm_6_6, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5[6]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_rsp_0,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_25_nl = MUX_v_6_2_2((SC_SRAM_CONFIG[14:9]),
      (rva_out_reg_data_15_9_sva_dfm_10[5:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl
      = MUX_v_6_2_2(6'b000000, PECore_DecodeAxiRead_switch_lp_mux_25_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_12_5_0 = MUX1HOT_v_6_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl,
      rva_out_reg_data_15_9_sva_dfm_6_5_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5[5:0]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_rsp_1,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_26_nl = MUX_v_2_2_2((SC_SRAM_CONFIG[21:20]),
      (rva_out_reg_data_23_17_sva_dfm_8[4:3]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl
      = MUX_v_2_2_2(2'b00, PECore_DecodeAxiRead_switch_lp_mux_26_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_14_4_3 = MUX1HOT_v_2_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl,
      rva_out_reg_data_23_17_sva_dfm_6_4_3, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5[4:3]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_1,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_27_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[19:17]),
      (rva_out_reg_data_23_17_sva_dfm_8[2:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl
      = MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_27_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_14_2_0 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl,
      rva_out_reg_data_23_17_sva_dfm_6_2_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5[2:0]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_2,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_20_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[30:28]),
      (rva_out_reg_data_30_25_sva_dfm_8[5:3]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl =
      MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_20_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_16_5_3 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl,
      rva_out_reg_data_30_25_sva_dfm_6_5_3, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5[5:3]),
      (weight_port_read_out_data_0_3_sva_dfm_5_rsp_0[2:0]), {PECore_PushAxiRsp_if_asn_79
      , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_28_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[27:25]),
      (rva_out_reg_data_30_25_sva_dfm_8[2:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl
      = MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_28_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_16_2_0 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl,
      rva_out_reg_data_30_25_sva_dfm_6_2_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5[2:0]),
      (weight_port_read_out_data_0_3_sva_dfm_5_rsp_1[3:1]), {PECore_PushAxiRsp_if_asn_79
      , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_131_nl
      = (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[94]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]));
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_132_nl
      = (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[94]) & (~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1_6
      = MUX_s_1_8_2(weight_port_read_out_data_0_2_sva_dfm_1_1_6, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1[6]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_131_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_132_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_141_nl
      = MUX_v_2_2_2(2'b00, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[93:92]), weight_mem_write_arbxbar_xbar_for_1_for_not_270_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_273_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_142_nl
      = MUX_v_2_2_2(2'b00, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[93:92]), weight_mem_write_arbxbar_xbar_for_1_for_not_273_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_s000000
      = MUX_v_2_8_2(weight_port_read_out_data_0_2_sva_dfm_1_1_5_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[5:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[5:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1[5:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1[5:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1[5:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_141_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_142_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_271_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_143_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[91:88]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_271_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_274_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_144_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[91:88]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_274_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_s000001
      = MUX_v_4_8_2(weight_port_read_out_data_0_2_sva_dfm_1_1_3_0, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_143_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_144_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign rva_out_reg_data_and_215_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_4_1_enexo;
  assign rva_out_reg_data_and_216_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_87_80_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_217_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_218_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_219_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_95_88_sva_dfm_4_2_3_enexo;
  assign rva_out_reg_data_and_220_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_119_112_sva_dfm_4_1_1_enexo;
  assign rva_out_reg_data_and_221_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_111_104_sva_dfm_4_1_1_enexo;
  assign rva_out_reg_data_and_222_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_223_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_1_1_enexo;
  assign and_695_ssc = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign nor_613_ssc = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign and_697_ssc = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  assign nor_614_ssc = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | weight_mem_run_3_for_land_3_lpi_1_dfm_2);
  assign and_699_ssc = weight_mem_run_3_for_land_2_lpi_1_dfm_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign nor_615_ssc = ~(weight_mem_run_3_for_land_2_lpi_1_dfm_2 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign rva_out_reg_data_119_112_sva_dfm_4_mx0w0_7 = MUX1HOT_s_1_3_2(rva_out_reg_data_119_112_sva_dfm_7_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[119]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_39_nl = MUX_v_7_2_2(7'b0000000, rva_out_reg_data_119_112_sva_dfm_6_6_0,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_119_112_sva_dfm_4_mx0w0_6_0 = MUX1HOT_v_7_3_2(while_if_while_if_and_39_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[118:112]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_111_104_sva_dfm_4_mx0w0_7 = MUX1HOT_s_1_3_2(rva_out_reg_data_111_104_sva_dfm_7_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[111]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_38_nl = MUX_v_7_2_2(7'b0000000, rva_out_reg_data_111_104_sva_dfm_6_6_0,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_111_104_sva_dfm_4_mx0w0_6_0 = MUX1HOT_v_7_3_2(while_if_while_if_and_38_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[110:104]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_87
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_87_80_sva_dfm_8_7 = rva_out_reg_data_87_80_sva_dfm_6_7
      & rva_in_reg_rw_sva_5;
  assign rva_out_reg_data_95_88_sva_dfm_8_7 = rva_out_reg_data_95_88_sva_dfm_6_7
      & rva_in_reg_rw_sva_5;
  assign rva_out_reg_data_95_88_sva_dfm_8_6 = rva_out_reg_data_95_88_sva_dfm_6_6
      & rva_in_reg_rw_sva_5;
  assign rva_out_reg_data_95_88_sva_dfm_8_5_4 = MUX_v_2_2_2(2'b00, rva_out_reg_data_95_88_sva_dfm_6_5_4,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_and_224_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_95_88_sva_dfm_4_1_3_enexo;
  assign rva_out_reg_data_and_225_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_119_112_sva_dfm_4_4_1_enexo;
  assign rva_out_reg_data_and_226_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_111_104_sva_dfm_4_4_1_enexo;
  assign rva_out_reg_data_and_227_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_228_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_103_96_sva_dfm_4_4_1_enexo;
  assign rva_out_reg_data_and_229_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_119_112_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_230_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_111_104_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_111_104_sva_dfm_7_7 = rva_out_reg_data_111_104_sva_dfm_6_7
      & rva_in_reg_rw_sva_5;
  assign rva_out_reg_data_119_112_sva_dfm_7_7 = rva_out_reg_data_119_112_sva_dfm_6_7
      & rva_in_reg_rw_sva_5;
  assign PECore_DecodeAxiRead_switch_lp_mux_19_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[23]),
      (rva_out_reg_data_23_17_sva_dfm_8[6]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl
      = PECore_DecodeAxiRead_switch_lp_mux_19_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_14_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl,
      rva_out_reg_data_23_17_sva_dfm_6_6, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5[6]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_0_1,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_29_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[22]),
      (rva_out_reg_data_23_17_sva_dfm_8[5]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_30_nl
      = PECore_DecodeAxiRead_switch_lp_mux_29_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_14_5 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_30_nl,
      rva_out_reg_data_23_17_sva_dfm_6_5, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5[5]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_0_0,
      {PECore_PushAxiRsp_if_asn_79 , PECore_PushAxiRsp_if_asn_81 , PECore_PushAxiRsp_if_asn_83
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign rva_out_reg_data_and_231_enex5 = rva_out_reg_data_and_25_cse & reg_rva_out_reg_data_95_88_sva_dfm_4_4_3_enexo;
  assign rva_out_reg_data_and_232_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_95_88_sva_dfm_4_3_3_enexo;
  assign or_dcpl_319 = weight_mem_run_3_for_5_and_143_itm_2 | weight_mem_run_3_for_5_and_142_itm_1;
  assign or_dcpl_323 = weight_mem_run_3_for_5_and_134_itm_2 | weight_mem_run_3_for_5_and_140_itm_2;
  assign or_dcpl_324 = weight_mem_run_3_for_5_and_136_itm_1 | weight_mem_run_3_for_5_and_135_itm_1;
  assign or_dcpl_332 = weight_mem_run_3_for_5_and_135_itm_1 | weight_mem_run_3_for_5_and_134_itm_2;
  assign or_dcpl_336 = weight_mem_run_3_for_5_and_142_itm_1 | weight_mem_run_3_for_5_and_140_itm_2;
  assign or_dcpl_337 = weight_mem_run_3_for_5_and_136_itm_1 | weight_mem_run_3_for_5_and_143_itm_2;
  assign or_tmp_586 = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  assign and_dcpl_886 = while_stage_0_3 & fsm_output;
  assign or_1125_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1;
  assign or_1124_nl = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1;
  assign mux_563_nl = MUX_s_1_2_2(or_1125_nl, or_1124_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign or_1123_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1;
  assign mux_564_nl = MUX_s_1_2_2(mux_563_nl, or_1123_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_tmp_622 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | mux_564_nl;
  assign or_tmp_623 = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | rva_in_reg_rw_sva_st_1_5 | (~ or_tmp_622);
  assign or_1128_cse = (~ while_stage_0_8) | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1;
  assign mux_565_cse = MUX_s_1_2_2(or_1128_cse, or_tmp_622, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign or_1141_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1;
  assign or_1140_nl = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1;
  assign mux_575_nl = MUX_s_1_2_2(or_1141_nl, or_1140_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign or_1139_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1;
  assign mux_576_nl = MUX_s_1_2_2(mux_575_nl, or_1139_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_tmp_638 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | mux_576_nl;
  assign or_tmp_639 = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | rva_in_reg_rw_sva_st_1_5 | (~ or_tmp_638);
  assign or_1144_nl = (~ while_stage_0_8) | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1;
  assign mux_577_itm = MUX_s_1_2_2(or_1144_nl, or_tmp_638, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_1641_cse = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
      | (~ while_stage_0_8) | weight_mem_run_3_for_land_1_lpi_1_dfm_3) & while_stage_0_7;
  assign and_1642_nl = or_1128_cse & while_stage_0_7;
  assign and_1643_nl = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1)
      & while_stage_0_7;
  assign and_1644_nl = ((~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1)
      & while_stage_0_7;
  assign mux_587_nl = MUX_s_1_2_2(and_1643_nl, and_1644_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign and_1645_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1)
      & while_stage_0_7;
  assign mux_588_nl = MUX_s_1_2_2(mux_587_nl, and_1645_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign mux_589_nl = MUX_s_1_2_2(and_1642_nl, mux_588_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign mux_tmp_546 = MUX_s_1_2_2(and_1641_cse, mux_589_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_1652_nl = ((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      | (~ while_stage_0_8) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1) & while_stage_0_7;
  assign and_1653_nl = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1)
      & while_stage_0_7;
  assign and_1654_nl = ((~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1)
      & while_stage_0_7;
  assign mux_601_nl = MUX_s_1_2_2(and_1653_nl, and_1654_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign and_1655_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1)
      & while_stage_0_7;
  assign mux_602_nl = MUX_s_1_2_2(mux_601_nl, and_1655_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign mux_603_nl = MUX_s_1_2_2(and_1652_nl, mux_602_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign mux_tmp_560 = MUX_s_1_2_2(and_1641_cse, mux_603_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_1657_nl = ((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6)
      | (~ while_stage_0_8) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1) & while_stage_0_7;
  assign and_1658_nl = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1)
      & while_stage_0_7;
  assign and_1659_nl = ((~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1)
      & while_stage_0_7;
  assign mux_608_nl = MUX_s_1_2_2(and_1658_nl, and_1659_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign and_1660_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1)
      & while_stage_0_7;
  assign mux_609_nl = MUX_s_1_2_2(mux_608_nl, and_1660_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign mux_610_nl = MUX_s_1_2_2(and_1657_nl, mux_609_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign mux_tmp_567 = MUX_s_1_2_2(and_1641_cse, mux_610_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign data_in_tmp_operator_2_for_and_tmp = PECoreRun_wen & weight_mem_run_3_for_land_2_lpi_1_dfm_2
      & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign data_in_tmp_operator_2_for_and_31_tmp = PECoreRun_wen & and_dcpl_33 & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign pe_manager_base_input_and_tmp = PECoreRun_wen & ((nand_88_cse & while_stage_0_3)
      | and_dcpl_220);
  assign rva_in_reg_data_and_tmp = PECoreRun_wen & and_dcpl_321 & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & (and_319_cse | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign input_mem_banks_read_1_read_data_and_4_tmp = PECoreRun_wen & (and_380_cse
      | ((~ reg_rva_in_reg_rw_sva_st_1_1_cse) & input_read_req_valid_lpi_1_dfm_1_1
      & and_dcpl_212));
  assign input_mem_banks_read_read_data_and_44_tmp = PECoreRun_wen & (~((~((~ rva_in_reg_rw_sva_st_1_4)
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)))
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
      & while_stage_0_6;
  assign or_1048_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (~((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:0]!=16'b0000000000000001)))
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ while_stage_0_3) | (~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1)));
  assign nor_638_nl = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])));
  assign mux_550_nl = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, or_1048_nl,
      nor_638_nl);
  assign and_1441_tmp = (~ mux_550_nl) & and_dcpl_220 & PECoreRun_wen;
  assign mux_579_nl = MUX_s_1_2_2((~ mux_577_itm), or_tmp_639, and_1624_cse);
  assign mux_578_nl = MUX_s_1_2_2((~ mux_577_itm), or_tmp_639, and_1625_cse);
  assign mux_580_nl = MUX_s_1_2_2(mux_579_nl, mux_578_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_1568_tmp = (~ mux_580_nl) & and_dcpl_41 & PECoreRun_wen;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_63_cse <= 1'b0;
      reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_56_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_act_port_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3
          <= 1'b0;
      pe_config_manager_counter_sva_dfm_3_1 <= 4'b0000;
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= 1'b0;
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= 1'b0;
      while_stage_0_3 <= 1'b0;
      while_stage_0_4 <= 1'b0;
      while_stage_0_5 <= 1'b0;
      while_stage_0_6 <= 1'b0;
      while_stage_0_7 <= 1'b0;
      while_stage_0_8 <= 1'b0;
      while_stage_0_9 <= 1'b0;
      while_stage_0_10 <= 1'b0;
      while_stage_0_11 <= 1'b0;
      while_stage_0_12 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1
          <= 1'b0;
      input_read_addrs_sva_1_1 <= 8'b00000000;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= 1'b0;
      weight_port_read_out_data_0_5_sva_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_4_sva_rsp_0 <= 1'b0;
      reg_weight_port_read_out_data_0_2_ftd <= 1'b0;
      reg_weight_port_read_out_data_0_2_ftd_1 <= 1'b0;
      weight_port_read_out_data_0_2_sva_5_4 <= 2'b00;
      weight_port_read_out_data_0_1_sva_7 <= 1'b0;
    end
    else if ( PECoreRun_wen ) begin
      reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_63_cse <= and_530_rmff;
      reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_56_cse <= and_533_rmff;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= and_537_rmff;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= and_541_rmff;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= and_545_rmff;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= and_549_rmff;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= and_554_rmff;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= and_558_rmff;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= and_563_rmff;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= and_566_rmff;
      reg_rva_out_Push_mioi_iswt0_cse <= and_568_cse;
      reg_start_PopNB_mioi_iswt0_cse <= and_570_rmff;
      reg_act_port_Push_mioi_iswt0_cse <= and_572_rmff;
      reg_rva_in_PopNB_mioi_iswt0_cse <= fsm_output;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_6
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_5
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_4
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
      pe_config_manager_counter_sva_dfm_3_1 <= MUX_v_4_2_2(4'b0000, operator_4_false_acc_nl,
          pe_config_UpdateManagerCounter_if_not_7_nl);
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= ~((pe_config_input_counter_sva_mx1 != (operator_16_false_acc_sdt_sva_1[7:0]))
          | (operator_16_false_acc_sdt_sva_1[8]));
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
      while_stage_0_3 <= reg_rva_in_PopNB_mioi_iswt0_cse;
      while_stage_0_4 <= while_stage_0_3;
      while_stage_0_5 <= while_stage_0_4;
      while_stage_0_6 <= while_stage_0_5;
      while_stage_0_7 <= while_stage_0_6;
      while_stage_0_8 <= while_stage_0_7;
      while_stage_0_9 <= while_stage_0_8;
      while_stage_0_10 <= while_stage_0_9;
      while_stage_0_11 <= while_stage_0_10;
      while_stage_0_12 <= while_stage_0_11;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1 <= ~ (pe_manager_base_weight_sva_mx2[1]);
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 <= pe_manager_base_weight_sva_mx3_0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1 <= pe_manager_base_weight_sva_mx2[1];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[2];
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= (pe_manager_base_weight_sva_mx1_3_0[2])
          & pe_manager_base_weight_sva_mx3_0 & (~ (pe_manager_base_weight_sva_mx2[1]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1
          <= ~((pe_manager_base_weight_sva_mx1_3_0[2]) | (pe_manager_base_weight_sva_mx2[1])
          | pe_manager_base_weight_sva_mx3_0);
      input_read_addrs_sva_1_1 <= nl_input_read_addrs_sva_1_1[7:0];
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
      weight_port_read_out_data_0_5_sva_rsp_0 <= weight_port_read_out_data_0_5_sva_mx0_7;
      weight_port_read_out_data_0_4_sva_rsp_0 <= weight_port_read_out_data_0_4_sva_mx0_7;
      reg_weight_port_read_out_data_0_2_ftd <= weight_port_read_out_data_0_2_sva_mx0_7;
      reg_weight_port_read_out_data_0_2_ftd_1 <= weight_port_read_out_data_0_2_sva_mx0_6;
      weight_port_read_out_data_0_2_sva_5_4 <= weight_port_read_out_data_0_2_sva_mx0_5_4;
      weight_port_read_out_data_0_1_sva_7 <= weight_port_read_out_data_0_1_sva_mx0_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_10 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_2_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_10 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_10 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_147_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_10 <= rva_out_reg_data_15_9_sva_dfm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_8 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_148_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_8 <= rva_out_reg_data_23_17_sva_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_8 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_149_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_8 <= rva_out_reg_data_30_25_sva_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_120_sva_dfm_4_5 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_150_enex5 ) begin
      rva_out_reg_data_127_120_sva_dfm_4_5 <= rva_out_reg_data_127_120_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_72_sva_dfm_4_5 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_151_enex5 ) begin
      rva_out_reg_data_79_72_sva_dfm_4_5 <= rva_out_reg_data_79_72_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_4_5 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_152_enex5 ) begin
      rva_out_reg_data_71_64_sva_dfm_4_5 <= rva_out_reg_data_71_64_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_63_sva_dfm_4_5 <= 1'b0;
      rva_out_reg_data_47_sva_dfm_4_5 <= 1'b0;
      input_read_req_valid_lpi_1_dfm_1_10 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_5_3 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_5_2_0 <= 3'b000;
      rva_out_reg_data_95_88_sva_dfm_4_5_rsp_0 <= 1'b0;
      rva_out_reg_data_87_80_sva_dfm_4_5_rsp_0 <= 1'b0;
      rva_out_reg_data_119_112_sva_dfm_4_5_rsp_0 <= 1'b0;
      rva_out_reg_data_111_104_sva_dfm_4_5_rsp_0 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_0 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_25_cse ) begin
      rva_out_reg_data_63_sva_dfm_4_5 <= rva_out_reg_data_63_sva_dfm_4_4;
      rva_out_reg_data_47_sva_dfm_4_5 <= rva_out_reg_data_47_sva_dfm_4_4;
      input_read_req_valid_lpi_1_dfm_1_10 <= input_read_req_valid_lpi_1_dfm_1_9;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
      rva_out_reg_data_39_36_sva_dfm_4_5_3 <= reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd;
      rva_out_reg_data_39_36_sva_dfm_4_5_2_0 <= reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1;
      rva_out_reg_data_95_88_sva_dfm_4_5_rsp_0 <= rva_out_reg_data_95_88_sva_dfm_4_4_7;
      rva_out_reg_data_87_80_sva_dfm_4_5_rsp_0 <= rva_out_reg_data_87_80_sva_dfm_4_4_7;
      rva_out_reg_data_119_112_sva_dfm_4_5_rsp_0 <= rva_out_reg_data_119_112_sva_dfm_4_4_7;
      rva_out_reg_data_111_104_sva_dfm_4_5_rsp_0 <= rva_out_reg_data_111_104_sva_dfm_4_4_7;
      rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_0 <= rva_out_reg_data_95_88_sva_dfm_4_4_6;
      rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_1 <= rva_out_reg_data_95_88_sva_dfm_4_4_5_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_153_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_5 <= rva_out_reg_data_62_56_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_5 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_154_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_5 <= rva_out_reg_data_35_32_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_5 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_155_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_5 <= rva_out_reg_data_55_48_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_156_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_5 <= rva_out_reg_data_46_40_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_6 <=
          1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_rsp_0
          <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_1
          <= 2'b00;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_2
          <= 3'b000;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_0_1
          <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_0_0
          <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_123_cse ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2 <= weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2 <= weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2 <= weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_6 <=
          reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_rsp_0
          <= weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_6;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_1
          <= weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_4_3;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_2
          <= weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_2_0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_0_1
          <= reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_rsp_0_0
          <= reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_47_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_48_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_49_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_50_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_10 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
          <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_cse ) begin
      rva_in_reg_rw_sva_10 <= rva_in_reg_rw_sva_9;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_10 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_4 ) begin
      rva_in_reg_rw_sva_st_1_10 <= rva_in_reg_rw_sva_st_1_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_8_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_16_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_31_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_24_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_7_1_sva_dfm_6_6 <= 1'b0;
      rva_out_reg_data_7_1_sva_dfm_6_5_0 <= 6'b000000;
      rva_out_reg_data_15_9_sva_dfm_6_6 <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_6_5_0 <= 6'b000000;
      rva_out_reg_data_23_17_sva_dfm_6_4_3 <= 2'b00;
      rva_out_reg_data_23_17_sva_dfm_6_2_0 <= 3'b000;
      rva_out_reg_data_30_25_sva_dfm_6_5_3 <= 3'b000;
      rva_out_reg_data_30_25_sva_dfm_6_2_0 <= 3'b000;
      rva_out_reg_data_23_17_sva_dfm_6_6 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_6_5 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_cse ) begin
      rva_out_reg_data_0_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_24_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
      rva_out_reg_data_8_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_25_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
      rva_out_reg_data_16_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_26_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
      rva_out_reg_data_31_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_17;
      rva_out_reg_data_24_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_15;
      rva_out_reg_data_7_1_sva_dfm_6_6 <= PECore_PushAxiRsp_if_mux1h_10_6;
      rva_out_reg_data_7_1_sva_dfm_6_5_0 <= PECore_PushAxiRsp_if_mux1h_10_5_0;
      rva_out_reg_data_15_9_sva_dfm_6_6 <= PECore_PushAxiRsp_if_mux1h_12_6;
      rva_out_reg_data_15_9_sva_dfm_6_5_0 <= PECore_PushAxiRsp_if_mux1h_12_5_0;
      rva_out_reg_data_23_17_sva_dfm_6_4_3 <= PECore_PushAxiRsp_if_mux1h_14_4_3;
      rva_out_reg_data_23_17_sva_dfm_6_2_0 <= PECore_PushAxiRsp_if_mux1h_14_2_0;
      rva_out_reg_data_30_25_sva_dfm_6_5_3 <= PECore_PushAxiRsp_if_mux1h_16_5_3;
      rva_out_reg_data_30_25_sva_dfm_6_2_0 <= PECore_PushAxiRsp_if_mux1h_16_2_0;
      rva_out_reg_data_23_17_sva_dfm_6_6 <= PECore_PushAxiRsp_if_mux1h_14_6;
      rva_out_reg_data_23_17_sva_dfm_6_5 <= PECore_PushAxiRsp_if_mux1h_14_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_16_0_sva_dfm_1_2 <= 17'b00000000000000000;
    end
    else if ( act_port_reg_data_and_19_enex5 ) begin
      act_port_reg_data_16_0_sva_dfm_1_2 <= act_port_reg_data_16_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_240_224_sva_dfm_1_2 <= 17'b00000000000000000;
    end
    else if ( act_port_reg_data_and_20_enex5 ) begin
      act_port_reg_data_240_224_sva_dfm_1_2 <= act_port_reg_data_240_224_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_48_32_sva_dfm_1_1 <= 17'b00000000000000000;
      act_port_reg_data_80_64_sva_dfm_1_1 <= 17'b00000000000000000;
      act_port_reg_data_112_96_sva_dfm_1_1 <= 17'b00000000000000000;
      act_port_reg_data_144_128_sva_dfm_1_1 <= 17'b00000000000000000;
    end
    else if ( and_1224_cse ) begin
      act_port_reg_data_48_32_sva_dfm_1_1 <= MUX_v_17_2_2((readslicef_28_17_11(PECore_RunScale_if_for_2_scaled_val_mul_1_nl)),
          act_port_reg_data_48_32_sva_mx1, or_dcpl_220);
      act_port_reg_data_80_64_sva_dfm_1_1 <= MUX_v_17_2_2((readslicef_28_17_11(PECore_RunScale_if_for_3_scaled_val_mul_1_nl)),
          act_port_reg_data_80_64_sva_mx1, or_dcpl_220);
      act_port_reg_data_112_96_sva_dfm_1_1 <= MUX_v_17_2_2((readslicef_28_17_11(PECore_RunScale_if_for_4_scaled_val_mul_1_nl)),
          act_port_reg_data_112_96_sva_mx1, or_dcpl_220);
      act_port_reg_data_144_128_sva_dfm_1_1 <= MUX_v_17_2_2((readslicef_28_17_11(PECore_RunScale_if_for_5_scaled_val_mul_1_nl)),
          act_port_reg_data_144_128_sva_mx1, or_dcpl_220);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_208_192_sva_dfm_1_2 <= 17'b00000000000000000;
    end
    else if ( act_port_reg_data_and_21_enex5 ) begin
      act_port_reg_data_208_192_sva_dfm_1_2 <= act_port_reg_data_208_192_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_176_160_sva_dfm_1_2 <= 17'b00000000000000000;
    end
    else if ( act_port_reg_data_and_22_enex5 ) begin
      act_port_reg_data_176_160_sva_dfm_1_2 <= act_port_reg_data_176_160_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_10 <= 1'b0;
    end
    else if ( PECore_PushOutput_if_and_cse ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_10 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_9 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_9 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= 1'b0;
      rva_in_reg_rw_sva_9 <= 1'b0;
    end
    else if ( while_if_and_6_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
      rva_in_reg_rw_sva_9 <= rva_in_reg_rw_sva_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_8 <= 1'b0;
      rva_in_reg_rw_sva_st_8 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_2_cse ) begin
      rva_in_reg_rw_sva_st_1_8 <= rva_in_reg_rw_sva_st_1_7;
      rva_in_reg_rw_sva_st_8 <= rva_in_reg_rw_sva_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_30 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_7)
        ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_1_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= 1'b0;
      rva_in_reg_rw_sva_8 <= 1'b0;
    end
    else if ( while_if_and_7_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
      rva_in_reg_rw_sva_8 <= rva_in_reg_rw_sva_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_2_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= 1'b0;
      weight_port_read_out_data_0_7_sva <= 8'b00000000;
      rva_in_reg_rw_sva_7 <= 1'b0;
      weight_port_read_out_data_0_5_sva_rsp_1 <= 7'b0000000;
      weight_port_read_out_data_0_4_sva_rsp_1 <= 7'b0000000;
      weight_port_read_out_data_0_3_sva_7_4 <= 4'b0000;
      weight_port_read_out_data_0_3_sva_3_0 <= 4'b0000;
      weight_port_read_out_data_0_2_sva_3_0 <= 4'b0000;
      weight_port_read_out_data_0_1_sva_6_0 <= 7'b0000000;
    end
    else if ( while_if_and_8_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6;
      weight_port_read_out_data_0_7_sva <= weight_port_read_out_data_0_7_sva_mx0;
      rva_in_reg_rw_sva_7 <= rva_in_reg_rw_sva_6;
      weight_port_read_out_data_0_5_sva_rsp_1 <= weight_port_read_out_data_0_5_sva_mx0_6_0;
      weight_port_read_out_data_0_4_sva_rsp_1 <= weight_port_read_out_data_0_4_sva_mx0_6_0;
      weight_port_read_out_data_0_3_sva_7_4 <= weight_port_read_out_data_0_3_sva_mx0_7_4;
      weight_port_read_out_data_0_3_sva_3_0 <= weight_port_read_out_data_0_3_sva_mx0_3_0;
      weight_port_read_out_data_0_2_sva_3_0 <= weight_port_read_out_data_0_2_sva_mx0_3_0;
      weight_port_read_out_data_0_1_sva_6_0 <= weight_port_read_out_data_0_1_sva_mx0_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_enex5 ) begin
      weight_port_read_out_data_1_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
          <= MUX_v_8_2_2(8'b00000000, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_2_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_3 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
          <= 1'b0;
      rva_in_reg_rw_sva_6 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_cse ) begin
      weight_mem_run_3_for_land_2_lpi_1_dfm_3 <= weight_mem_run_3_for_land_2_lpi_1_dfm_2;
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= weight_mem_run_3_for_land_3_lpi_1_dfm_2;
      weight_mem_run_3_for_land_5_lpi_1_dfm_3 <= weight_mem_run_3_for_land_5_lpi_1_dfm_2;
      weight_mem_run_3_for_land_4_lpi_1_dfm_3 <= weight_mem_run_3_for_land_4_lpi_1_dfm_2;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_6
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
      rva_in_reg_rw_sva_6 <= rva_in_reg_rw_sva_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_190_enex5 ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_191_enex5 ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_192_enex5 ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_3_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_193_enex5 ) begin
      weight_port_read_out_data_2_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_4_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_194_enex5 ) begin
      weight_port_read_out_data_2_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_5_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_195_enex5 ) begin
      weight_port_read_out_data_2_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_196_enex5 ) begin
      weight_port_read_out_data_2_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_7_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_197_enex5 ) begin
      weight_port_read_out_data_2_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_8_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_198_enex5 ) begin
      weight_port_read_out_data_2_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_9_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_199_enex5 ) begin
      weight_port_read_out_data_2_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_10_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_200_enex5 ) begin
      weight_port_read_out_data_2_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_11_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_201_enex5 ) begin
      weight_port_read_out_data_2_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_12_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_202_enex5 ) begin
      weight_port_read_out_data_2_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_13_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_203_enex5 ) begin
      weight_port_read_out_data_2_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_204_enex5 ) begin
      weight_port_read_out_data_2_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_205_enex5 ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
          <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[7:0]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[15:8]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[23:16]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[31:24]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[39:32]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[47:40]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[55:48]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[71:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[71:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[71:64]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[71:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[63:56]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:72]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:72]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:72]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:72]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[71:64]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[87:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[87:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[87:80]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[87:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[79:72]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:88]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:88]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:88]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:88]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[87:80]),
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[103:96]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[103:96]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[103:96]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[103:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[103:96]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[95:88]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:104]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:104]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:104]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:104]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:104]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[103:96]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[119:112]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[119:112]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[119:112]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[119:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[119:112]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[111:104]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_206_enex5 ) begin
      weight_port_read_out_data_4_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_2_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_207_enex5 ) begin
      weight_port_read_out_data_4_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_3_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_208_enex5 ) begin
      weight_port_read_out_data_4_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_4_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_209_enex5 ) begin
      weight_port_read_out_data_4_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_5_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_210_enex5 ) begin
      weight_port_read_out_data_4_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_211_enex5 ) begin
      weight_port_read_out_data_4_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_7_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_212_enex5 ) begin
      weight_port_read_out_data_4_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_8_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_213_enex5 ) begin
      weight_port_read_out_data_4_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_9_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_214_enex5 ) begin
      weight_port_read_out_data_4_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_10_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_215_enex5 ) begin
      weight_port_read_out_data_4_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_11_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_216_enex5 ) begin
      weight_port_read_out_data_4_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_12_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_217_enex5 ) begin
      weight_port_read_out_data_4_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_13_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_218_enex5 ) begin
      weight_port_read_out_data_4_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_219_enex5 ) begin
      weight_port_read_out_data_4_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_31_enex5 ) begin
      weight_port_read_out_data_3_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_31_tmp ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000
          <= MUX_v_8_2_2(8'b00000000, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_1_nl,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_3_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_5,
          (weight_port_read_out_data_0_7_sva_dfm_mx0w2[7]), PECore_PushAxiRsp_if_else_mux_23_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_40_tmp , while_and_39_cse});
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5,
          weight_port_read_out_data_0_5_sva_dfm_mx0w2_7, PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_40_tmp , while_and_39_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        & while_stage_0_6 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        & while_stage_0_6 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_5 <= 1'b0;
      rva_in_reg_rw_sva_st_5 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_3_cse ) begin
      rva_in_reg_rw_sva_st_1_5 <= rva_in_reg_rw_sva_st_1_4;
      rva_in_reg_rw_sva_st_5 <= rva_in_reg_rw_sva_st_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2 <= 1'b0;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_140_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_142_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_143_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_134_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_135_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_136_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_100_itm_1 <= 1'b0;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= 3'b000;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_12_itm_1 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_14_itm_1_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_15_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_16_itm_1_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_4_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_6_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_7_itm_1 <= 1'b0;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_146_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_147_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_148_itm_2 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_149_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_2 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_151_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_152_itm_2_cse <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= 1'b0;
    end
    else if ( weight_mem_banks_read_1_read_data_and_8_cse ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_140_itm_2 <= weight_mem_run_3_for_5_and_140_itm_1;
      weight_mem_run_3_for_5_and_142_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_143_itm_2 <= weight_mem_run_3_for_5_and_143_itm_1;
      weight_mem_run_3_for_5_and_134_itm_2 <= weight_mem_run_3_for_5_and_134_itm_1;
      weight_mem_run_3_for_5_and_135_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_136_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b111)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_15_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_2_2_0!=3'b000));
      weight_mem_run_3_for_5_and_100_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b011)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= weight_read_addrs_7_lpi_1_dfm_2_2_0;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
      weight_mem_run_3_for_5_and_12_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1;
      reg_weight_mem_run_3_for_5_and_14_itm_1_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1;
      reg_weight_mem_run_3_for_5_and_15_itm_2_cse <= weight_mem_run_3_for_5_and_15_itm_1;
      reg_weight_mem_run_3_for_5_and_16_itm_1_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1;
      reg_weight_mem_run_3_for_5_and_4_itm_2_cse <= weight_mem_run_3_for_5_and_4_itm_1;
      reg_weight_mem_run_3_for_5_and_6_itm_2_cse <= weight_mem_run_3_for_5_and_6_itm_1;
      weight_mem_run_3_for_5_and_7_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_2_cse <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1;
      reg_weight_mem_run_3_for_5_and_146_itm_2_cse <= weight_mem_run_3_for_5_and_146_itm_1;
      reg_weight_mem_run_3_for_5_and_147_itm_2_cse <= weight_mem_run_3_for_5_and_147_itm_1;
      weight_mem_run_3_for_5_and_148_itm_2 <= weight_mem_run_3_for_5_and_148_itm_1;
      reg_weight_mem_run_3_for_5_and_149_itm_2_cse <= weight_mem_run_3_for_5_and_149_itm_1;
      weight_mem_run_3_for_5_and_150_itm_2 <= weight_mem_run_3_for_5_and_150_itm_1;
      reg_weight_mem_run_3_for_5_and_151_itm_2_cse <= weight_mem_run_3_for_5_and_151_itm_1;
      reg_weight_mem_run_3_for_5_and_152_itm_2_cse <= weight_mem_run_3_for_5_and_152_itm_1;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= weight_read_addrs_5_lpi_1_dfm_2_2_0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & weight_mem_run_3_for_land_7_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_7_nl & while_stage_0_6 ) begin
      reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2_cse <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_1_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_6_sva_dfm_2 <= 8'b00000000;
      weight_port_read_out_data_0_8_sva_dfm_2 <= 8'b00000000;
      weight_port_read_out_data_0_9_sva_dfm_2 <= 8'b00000000;
      weight_port_read_out_data_0_15_sva_dfm_2 <= 8'b00000000;
      weight_port_read_out_data_0_10_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_10_sva_dfm_2_6_0 <= 7'b0000000;
      weight_port_read_out_data_0_11_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_11_sva_dfm_2_6 <= 1'b0;
      weight_port_read_out_data_0_11_sva_dfm_2_5_4 <= 2'b00;
      weight_port_read_out_data_0_11_sva_dfm_2_3_0 <= 4'b0000;
      weight_port_read_out_data_0_12_sva_dfm_2_7_4 <= 4'b0000;
      weight_port_read_out_data_0_12_sva_dfm_2_3_0 <= 4'b0000;
      weight_port_read_out_data_0_13_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_13_sva_dfm_2_6_0 <= 7'b0000000;
      weight_port_read_out_data_0_14_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_14_sva_dfm_2_6_0 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_136_cse ) begin
      weight_port_read_out_data_0_6_sva_dfm_2 <= MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_sva_1,
          while_and_40_tmp);
      weight_port_read_out_data_0_8_sva_dfm_2 <= MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_63_56_sva_1,
          while_and_40_tmp);
      weight_port_read_out_data_0_9_sva_dfm_2 <= MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_71_64_sva_1,
          while_and_40_tmp);
      weight_port_read_out_data_0_15_sva_dfm_2 <= MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_119_112_sva_1,
          while_and_40_tmp);
      weight_port_read_out_data_0_10_sva_dfm_2_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010[7]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_sva_1_7,
          while_and_40_tmp);
      weight_port_read_out_data_0_10_sva_dfm_2_6_0 <= MUX_v_7_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010[6:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_79_72_s000000,
          while_and_40_tmp);
      weight_port_read_out_data_0_11_sva_dfm_2_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009[7]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1_7,
          while_and_40_tmp);
      weight_port_read_out_data_0_11_sva_dfm_2_6 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009[6]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_sva_1_6,
          while_and_40_tmp);
      weight_port_read_out_data_0_11_sva_dfm_2_5_4 <= MUX_v_2_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009[5:4]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_s000000,
          while_and_40_tmp);
      weight_port_read_out_data_0_11_sva_dfm_2_3_0 <= MUX_v_4_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009[3:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_87_80_s000001,
          while_and_40_tmp);
      weight_port_read_out_data_0_12_sva_dfm_2_7_4 <= MUX_v_4_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012[7:4]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_s000000,
          while_and_40_tmp);
      weight_port_read_out_data_0_12_sva_dfm_2_3_0 <= MUX_v_4_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012[3:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_95_88_s000001,
          while_and_40_tmp);
      weight_port_read_out_data_0_13_sva_dfm_2_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011[7]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000000,
          while_and_40_tmp);
      weight_port_read_out_data_0_13_sva_dfm_2_6_0 <= MUX_v_7_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011[6:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_103_96_000001,
          while_and_40_tmp);
      weight_port_read_out_data_0_14_sva_dfm_2_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014[7]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000000,
          while_and_40_tmp);
      weight_port_read_out_data_0_14_sva_dfm_2_6_0 <= MUX_v_7_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014[6:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_111_104000001,
          while_and_40_tmp);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= 1'b0;
      rva_in_reg_rw_sva_5 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_4_cse ) begin
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= weight_mem_run_3_for_land_1_lpi_1_dfm_2;
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= weight_mem_run_3_for_land_7_lpi_1_dfm_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= weight_mem_run_3_for_land_3_lpi_1_dfm_1;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= weight_mem_run_3_for_land_5_lpi_1_dfm_1;
      rva_in_reg_rw_sva_5 <= rva_in_reg_rw_sva_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_9_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_10_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_11_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_12_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_13_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_14_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_41_cse ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_nc000000;
      weight_port_read_out_data_6_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
      weight_port_read_out_data_6_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_n000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_9_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_10_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_11_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_12_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_13_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_145_cse ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
      weight_port_read_out_data_1_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
      weight_port_read_out_data_1_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
      weight_port_read_out_data_1_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
      weight_port_read_out_data_1_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
      weight_port_read_out_data_1_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
      weight_port_read_out_data_1_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
      weight_port_read_out_data_1_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
      weight_port_read_out_data_1_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
      weight_port_read_out_data_1_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
      weight_port_read_out_data_1_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
      weight_port_read_out_data_1_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
      weight_port_read_out_data_1_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
      weight_port_read_out_data_1_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
      weight_port_read_out_data_1_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_9_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_10_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_11_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_12_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_13_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_159_cse ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
      weight_port_read_out_data_5_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
      weight_port_read_out_data_5_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
      weight_port_read_out_data_5_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
      weight_port_read_out_data_5_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
      weight_port_read_out_data_5_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
      weight_port_read_out_data_5_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
      weight_port_read_out_data_5_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
      weight_port_read_out_data_5_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
      weight_port_read_out_data_5_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
      weight_port_read_out_data_5_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
      weight_port_read_out_data_5_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
      weight_port_read_out_data_5_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
      weight_port_read_out_data_5_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_9_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_10_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_11_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_12_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_13_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_85_cse ) begin
      weight_port_read_out_data_3_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001;
      weight_port_read_out_data_3_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000;
      weight_port_read_out_data_3_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003;
      weight_port_read_out_data_3_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002;
      weight_port_read_out_data_3_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005;
      weight_port_read_out_data_3_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004;
      weight_port_read_out_data_3_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000007;
      weight_port_read_out_data_3_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000006;
      weight_port_read_out_data_3_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000009;
      weight_port_read_out_data_3_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000008;
      weight_port_read_out_data_3_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000011;
      weight_port_read_out_data_3_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000010;
      weight_port_read_out_data_3_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000013;
      weight_port_read_out_data_3_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000012;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1244_cse | or_dcpl_319 | weight_mem_run_3_for_5_and_140_itm_2)
        & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_15_sva_dfm_1 <= weight_port_read_out_data_7_15_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1249_cse | or_dcpl_324 | or_dcpl_323) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_14_sva_dfm_1 <= weight_port_read_out_data_7_14_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_13_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1254_cse | weight_mem_run_3_for_5_and_135_itm_1 | weight_mem_run_3_for_5_and_142_itm_1
        | weight_mem_run_3_for_5_and_140_itm_2) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_13_sva_dfm_1 <= weight_port_read_out_data_7_13_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_12_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1254_cse | or_dcpl_332 | weight_mem_run_3_for_5_and_140_itm_2)
        & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_12_sva_dfm_1 <= weight_port_read_out_data_7_12_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_11_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1249_cse | or_dcpl_337 | or_dcpl_336) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_11_sva_dfm_1 <= weight_port_read_out_data_7_11_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_10_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1249_cse | or_dcpl_324 | weight_mem_run_3_for_5_and_134_itm_2
        | weight_mem_run_3_for_5_and_100_itm_1) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_10_sva_dfm_1 <= weight_port_read_out_data_7_10_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_9_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1274_cse | or_dcpl_324 | or_dcpl_336) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_9_sva_dfm_1 <= weight_port_read_out_data_7_9_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_8_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1280_cse ) begin
      weight_port_read_out_data_7_8_sva_dfm_1 <= weight_port_read_out_data_7_8_sva_dfm_3;
      weight_port_read_out_data_7_1_sva_dfm_1 <= weight_port_read_out_data_7_1_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_4_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1285_cse ) begin
      weight_port_read_out_data_7_7_sva_dfm_1 <= weight_port_read_out_data_7_7_sva_dfm_3;
      weight_port_read_out_data_7_6_sva_dfm_1 <= weight_port_read_out_data_7_6_sva_dfm_3;
      weight_port_read_out_data_7_5_sva_dfm_1 <= weight_port_read_out_data_7_5_sva_dfm_3;
      weight_port_read_out_data_7_4_sva_dfm_1 <= weight_port_read_out_data_7_4_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_3_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1254_cse | or_dcpl_332 | weight_mem_run_3_for_5_and_100_itm_1)
        & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_3_sva_dfm_1 <= weight_port_read_out_data_7_3_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_2_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1254_cse | or_dcpl_319 | weight_mem_run_3_for_5_and_100_itm_1)
        & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_2_sva_dfm_1 <= weight_port_read_out_data_7_2_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1274_cse | or_dcpl_324 | weight_mem_run_3_for_5_and_142_itm_1
        | weight_mem_run_3_for_5_and_100_itm_1) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_7_0_sva_dfm_1 <= weight_port_read_out_data_7_0_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1324_cse | reg_weight_mem_run_3_for_5_and_16_itm_1_cse | reg_weight_mem_run_3_for_5_and_15_itm_2_cse
        | reg_weight_mem_run_3_for_5_and_14_itm_1_cse | weight_mem_run_3_for_5_and_12_itm_1)
        & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_5_15_sva_dfm_1 <= weight_port_read_out_data_5_15_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1324_cse | reg_weight_mem_run_3_for_5_and_16_itm_1_cse | weight_mem_run_3_for_5_and_7_itm_1
        | reg_weight_mem_run_3_for_5_and_6_itm_2_cse | reg_weight_mem_run_3_for_5_and_4_itm_2_cse)
        & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_5_14_sva_dfm_1 <= weight_port_read_out_data_5_14_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_44_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_44_itm_1
          <= ~((weight_read_addrs_5_lpi_1_dfm_2_2_0!=3'b000));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_372_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_300_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_302_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2
          <= MUX_s_1_2_2(weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_10_nl & while_stage_0_6 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
          <= 1'b0;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_380_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
          <= ~((weight_read_addrs_3_lpi_1_dfm_2_2_0!=3'b000));
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= weight_read_addrs_3_lpi_1_dfm_2_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_384_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_136_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_134_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_151_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_2
          <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_389_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_1
          <= crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 <= 1'b0;
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_390_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_28_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_2 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_2 <= 1'b0;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2_cse <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_118_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_1;
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_2_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= 8'b00000000;
    end
    else if ( mux_539_nl & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_11_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= MUX_v_8_2_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[7:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_48_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_12_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= MUX_v_8_2_2((weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[7:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_80_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_8 <= 120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_231 | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & mux_18_nl ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_8 <= weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:8];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_231 | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & mux_24_nl ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_RunFSM_switch_lp_equal_tmp_1_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_UpdateFSM_switch_lp_equal_tmp_2_3 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_empty_sva_1[2])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_25_nl) & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_28_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1 <= 1'b0;
    end
    else if ( weight_read_addrs_and_5_cse ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_83 & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= 1'b0;
      rva_in_reg_rw_sva_4 <= 1'b0;
    end
    else if ( while_if_and_11_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp |
          Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp |
          Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_1
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_1
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_1
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_1
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= weight_mem_run_3_for_weight_mem_run_3_for_and_1_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_1
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= weight_mem_run_3_for_weight_mem_run_3_for_and_6_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_1
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0_1 | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & weight_mem_read_arbxbar_xbar_1_for_3_8_for_3_or_cse;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse;
      rva_in_reg_rw_sva_4 <= rva_in_reg_rw_sva_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_49_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_55_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_61_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_67_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse & (and_dcpl_83 | Arbiter_8U_Roundrobin_pick_and_25_cse)
        & or_dcpl_80 ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0,
          Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1, Arbiter_8U_Roundrobin_pick_and_25_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_73_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_78_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_84_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_90_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva <= 15'b000000000000000;
    end
    else if ( (~ mux_541_nl) & fsm_output & while_stage_0_5 & PECoreRun_wen ) begin
      pe_manager_base_weight_sva <= pe_manager_base_weight_sva_mx2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= 11'b00000000000;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= 1'b0;
    end
    else if ( weight_read_addrs_and_7_cse ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= MUX_v_11_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl,
          weight_read_addrs_0_14_4_lpi_1_dfm_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= MUX_s_1_2_2((weight_read_addrs_0_3_0_lpi_1_dfm_4[3]),
          (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_172 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_172 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_48_enex5 ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_15_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_49_enex5 ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_14_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_50_enex5 ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_13_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_51_enex5 ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_12_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_52_enex5 ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_11_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_53_enex5 ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_10_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_54_enex5 ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_9_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_55_enex5 ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_8_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_56_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_57_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_58_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_59_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_60_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_61_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_62_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_63_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= 12'b000000000000;
    end
    else if ( weight_write_addrs_and_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= weight_write_addrs_lpi_1_dfm_1_2[14:3];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= 1'b0;
      weight_read_addrs_1_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_3_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= 13'b0000000000000;
      weight_read_addrs_5_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_7_lpi_1_dfm_1 <= 15'b000000000000000;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1,
          and_162_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1,
          and_162_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1,
          and_162_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1,
          and_162_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1,
          and_162_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1,
          and_162_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1,
          and_162_cse);
      weight_read_addrs_1_lpi_1_dfm_1 <= weight_read_addrs_1_lpi_1_dfm_1_1;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_3_lpi_1_dfm_1 <= weight_read_addrs_3_lpi_1_dfm_1_1;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_1 <= weight_read_addrs_5_lpi_1_dfm_1_1;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_7_lpi_1_dfm_1 <= weight_read_addrs_7_lpi_1_dfm_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_15_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_not_185,
          weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0, and_113_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0, and_120_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0, and_127_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0, and_134_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0, and_141_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0, and_148_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0, and_dcpl_643);
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0, and_162_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1 <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= 1'b0;
      rva_in_reg_rw_sva_3 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= 1'b0;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1 <= MUX_s_1_2_2((pe_manager_base_weight_sva_mx1_3_0[2]),
          reg_rva_in_reg_rw_sva_2_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      rva_in_reg_rw_sva_3 <= reg_rva_in_reg_rw_sva_2_cse;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_55_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= 1'b0;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= 8'b00000000;
      rva_in_reg_rw_sva_st_3 <= 1'b0;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_1_for_and_cse ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_55_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b101)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b011)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b110)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= weight_mem_write_arbxbar_xbar_for_lshift_tmp;
      rva_in_reg_rw_sva_st_3 <= reg_rva_in_reg_rw_sva_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_and_cse ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_600);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_600);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_600);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_600);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_600);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_600);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_600);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_600);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_50_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_64_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse & ((~ while_stage_0_5) | while_and_1263_itm_1)
        ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= MUX_v_15_2_2(pe_manager_base_weight_sva_mx2,
          PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1, while_and_1263_itm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_64_enex5 ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_15_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_65_enex5 ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_14_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_66_enex5 ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_13_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_67_enex5 ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_12_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_68_enex5 ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_11_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_69_enex5 ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_10_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_70_enex5 ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_9_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_71_enex5 ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_8_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_72_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_7_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_73_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_6_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_74_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_5_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_75_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_76_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_3_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_77_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_2_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_78_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_1_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_79_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= 15'b000000000000000;
    end
    else if ( weight_write_addrs_and_2_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= pe_manager_base_input_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( weight_write_data_data_and_16_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_2_cse <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= 1'b0;
      while_and_1263_itm_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_4_cse ) begin
      reg_rva_in_reg_rw_sva_2_cse <= reg_rva_in_reg_rw_sva_st_1_1_cse;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= MUX_s_1_2_2(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
      while_and_1263_itm_1 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1
          & PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
          & reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= 4'b0000;
    end
    else if ( weight_read_addrs_and_29_enex5 ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= 11'b00000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_216 ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_2_1_sva <= 2'b00;
      pe_config_is_zero_first_sva <= 1'b0;
    end
    else if ( state_and_cse ) begin
      state_2_1_sva <= state_mux_1_cse;
      pe_config_is_zero_first_sva <= pe_config_is_zero_first_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_0_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_237) ) begin
      state_0_sva <= PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_manager_counter_sva <= 4'b0000;
    end
    else if ( (((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4:2]!=3'b000))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:5]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10:8]!=3'b000))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:11]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
        & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])
        & rva_in_PopNB_mioi_return_rsc_z_mxwt & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]))
        & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))
        & reg_rva_in_PopNB_mioi_iswt0_cse) | and_1341_cse) & PECoreRun_wen ) begin
      pe_config_manager_counter_sva <= MUX_v_4_2_2(pe_config_manager_counter_sva_dfm_3_1,
          PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl,
          and_662_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_num_manager_sva <= 4'b0001;
      pe_config_num_output_sva <= 8'b00000001;
    end
    else if ( pe_config_num_manager_and_cse ) begin
      pe_config_num_manager_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[35:32];
      pe_config_num_output_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= 1'b0;
      state_2_1_sva_dfm_1 <= 2'b00;
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= 8'b00000000;
      input_write_req_valid_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_5_cse ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= rva_in_PopNB_mioi_return_rsc_z_mxwt;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
      state_2_1_sva_dfm_1 <= MUX_v_2_2_2(PECore_UpdateFSM_switch_lp_and_1_nl, state_mux_1_cse,
          rva_in_PopNB_mioi_return_rsc_z_mxwt);
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= and_319_cse;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0];
      input_write_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= 1'b0;
      PECore_RunFSM_switch_lp_nor_tmp_1 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_9_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= PECore_UpdateFSM_switch_lp_equal_tmp_6;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= ~(PECore_RunScale_PECore_RunScale_if_and_1_svs_1
          | PECore_UpdateFSM_switch_lp_nor_tmp_1);
      PECore_RunFSM_switch_lp_nor_tmp_1 <= ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
          | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(or_380_cse | or_dcpl_237)) ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= input_port_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva <= 8'b00000000;
    end
    else if ( ((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
        | (~ reg_rva_in_PopNB_mioi_iswt0_cse) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
        | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)) & mux_542_nl & and_dcpl_886 &
        PECoreRun_wen ) begin
      pe_config_input_counter_sva <= pe_config_input_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva <= 8'b00000000;
    end
    else if ( (~((~((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
        | (~ reg_rva_in_PopNB_mioi_iswt0_cse) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
        | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt))) | mux_543_nl)) & and_dcpl_886
        & PECoreRun_wen ) begin
      pe_config_output_counter_sva <= pe_config_output_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      operator_8_false_acc_sdt_sva_1 <= 9'b000000000;
    end
    else if ( pe_config_UpdateManagerCounter_if_if_and_enex5 ) begin
      operator_8_false_acc_sdt_sva_1 <= nl_operator_8_false_acc_sdt_sva_1[8:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiWrite_switch_lp_and_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_48_32_sva <= 17'b00000000000000000;
      act_port_reg_data_80_64_sva <= 17'b00000000000000000;
      act_port_reg_data_112_96_sva <= 17'b00000000000000000;
      act_port_reg_data_144_128_sva <= 17'b00000000000000000;
    end
    else if ( and_1374_cse ) begin
      act_port_reg_data_48_32_sva <= act_port_reg_data_48_32_sva_mx1;
      act_port_reg_data_80_64_sva <= act_port_reg_data_80_64_sva_mx1;
      act_port_reg_data_112_96_sva <= act_port_reg_data_112_96_sva_mx1;
      act_port_reg_data_144_128_sva <= act_port_reg_data_144_128_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_1_19_0_sva <= 20'b00000000000000000000;
      accum_vector_data_2_19_0_sva <= 20'b00000000000000000000;
      accum_vector_data_4_19_0_sva <= 20'b00000000000000000000;
      accum_vector_data_3_19_0_sva <= 20'b00000000000000000000;
    end
    else if ( and_1393_cse ) begin
      accum_vector_data_1_19_0_sva <= MUX_v_20_2_2(20'b00000000000000000000, ProductSum_for_acc_38_nl,
          PECore_UpdateFSM_switch_lp_not_21_nl);
      accum_vector_data_2_19_0_sva <= MUX_v_20_2_2(20'b00000000000000000000, ProductSum_for_acc_30_nl,
          PECore_UpdateFSM_switch_lp_not_36_nl);
      accum_vector_data_4_19_0_sva <= MUX_v_20_2_2(20'b00000000000000000000, ProductSum_for_acc_26_nl,
          PECore_UpdateFSM_switch_lp_not_34_nl);
      accum_vector_data_3_19_0_sva <= MUX_v_20_2_2(20'b00000000000000000000, ProductSum_for_acc_22_nl,
          PECore_UpdateFSM_switch_lp_not_35_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0
          <= 7'b0000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( and_1415_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1
          <= MUX1HOT_v_8_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000005,
          weight_port_read_out_data_0_7_sva_mx0, {and_dcpl_583 , and_dcpl_655 , and_dcpl_656});
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_6_0
          <= MUX1HOT_v_7_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_138_nl,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003[6:0]),
          weight_port_read_out_data_0_5_sva_mx0_6_0, {and_dcpl_583 , and_dcpl_655
          , and_dcpl_656});
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_6_0
          <= MUX1HOT_v_7_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_137_nl,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004[6:0]),
          weight_port_read_out_data_0_4_sva_mx0_6_0, {and_dcpl_583 , and_dcpl_655
          , and_dcpl_656});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_1_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_249_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_174_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_189_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_204_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[127:120]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_219_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_250_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_175_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_190_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_205_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[119:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_220_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_251_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_176_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_191_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_206_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[111:104]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_221_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_252_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_177_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_192_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_207_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[103:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_222_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_253_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_178_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_193_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_208_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[95:88]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_223_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_254_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_179_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_194_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_209_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[87:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_224_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_240_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_255_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_180_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_195_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_210_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_225_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_241_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_181_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_196_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_211_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[79:72]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_226_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_242_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_257_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_182_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_197_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_212_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[71:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_227_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_51_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_243_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_244_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_246_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~ mux_tmp_31) & and_dcpl_48 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
        ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= MUX_v_8_2_2(8'b00000000, mux1h_3_nl, not_2374_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_53_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_198_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_201_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[23:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_202_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[15:8]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_203_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_54_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_228_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_229_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_231_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[15:8]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_233_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_57_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_199_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_200_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_59_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_245_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[7:0]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_140_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_62_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_230_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[23:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_232_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= 1'b0;
    end
    else if ( weight_read_addrs_and_17_cse ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= 1'b0;
    end
    else if ( PECoreRun_wen & weight_mem_run_3_for_land_5_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2 <= 2'b00;
    end
    else if ( PECoreRun_wen & mux_42_nl & while_stage_0_6 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2 <= MUX_v_2_2_2(pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_2[7:6]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_231 | (~ weight_mem_run_3_for_land_3_lpi_1_dfm_2)))
        ) begin
      weight_port_read_out_data_2_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_15_sva_dfm_1 <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_231 | (~ weight_mem_run_3_for_land_5_lpi_1_dfm_2)))
        ) begin
      weight_port_read_out_data_4_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_14_sva_dfm_1 <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_233 | (~ fsm_output))) & ((~ weight_mem_run_3_for_land_4_lpi_1_dfm_1)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        | (~ while_stage_0_6)) ) begin
      weight_port_read_out_data_3_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_5_and_143_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_140_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_134_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_15_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_6_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_4_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_152_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_151_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_149_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_148_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_147_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_146_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= 1'b0;
    end
    else if ( weight_read_addrs_and_19_cse ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= weight_read_addrs_7_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= weight_mem_run_3_for_weight_mem_run_3_for_and_7_tmp;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= weight_read_addrs_5_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_5_and_143_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b110)
          & weight_mem_run_3_for_weight_mem_run_3_for_and_7_tmp;
      weight_mem_run_3_for_5_and_140_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_weight_mem_run_3_for_and_7_tmp;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_134_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b101)
          & weight_mem_run_3_for_weight_mem_run_3_for_and_7_tmp;
      weight_mem_run_3_for_5_and_15_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= ~((weight_read_addrs_5_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_6_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1;
      weight_mem_run_3_for_5_and_4_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1_1;
      weight_mem_run_3_for_5_and_152_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
      weight_mem_run_3_for_5_and_151_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1;
      weight_mem_run_3_for_5_and_150_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1
          & (pe_manager_base_weight_sva[1:0]==2'b01) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_149_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
      weight_mem_run_3_for_5_and_148_itm_1 <= (pe_manager_base_weight_sva[1]) & PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          & (~ (pe_manager_base_weight_sva[2])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_147_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
      weight_mem_run_3_for_5_and_146_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1 <= ~((pe_manager_base_weight_sva[2:0]!=3'b000));
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_1
          <= 1'b0;
    end
    else if ( weight_read_addrs_and_21_cse ) begin
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= weight_read_addrs_3_lpi_1_dfm_1[2:0];
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_1
          <= ~((weight_read_addrs_3_lpi_1_dfm_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_43_nl ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_44_nl ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_61_nl ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_80_nl ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_89_nl ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_93_nl ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_30_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= 1'b0;
    end
    else if ( operator_15_false_1_and_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_162_cse | or_dcpl_75)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_dcpl_643 | or_dcpl_75)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_148_cse | or_dcpl_75)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_141_cse | or_dcpl_75)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_134_cse | or_dcpl_75)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_127_cse | or_dcpl_75)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_120_cse | or_dcpl_75)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= 15'b000000000000000;
    end
    else if ( PEManager_15U_PEManagerWrite_and_enex5 ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= rva_in_reg_data_sva_1[30:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_num_input_sva <= 8'b00000001;
      pe_manager_base_bias_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_num_input_and_cse ) begin
      pe_manager_num_input_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      pe_manager_base_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[46:32];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_is_valid_sva <= 1'b0;
      pe_config_is_cluster_sva <= 1'b0;
      pe_config_is_bias_sva <= 1'b0;
    end
    else if ( pe_config_is_valid_and_cse ) begin
      pe_config_is_valid_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
      pe_config_is_cluster_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[16];
      pe_config_is_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_zero_active_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & and_319_cse & (~ PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)
        & (~ or_dcpl_256) ) begin
      pe_manager_zero_active_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:2]==8'b00000000) & nor_721_cse
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:12]!=2'b00))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:14]!=2'b00)))
        & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]))
        | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
        | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 | (~(reg_rva_in_reg_rw_sva_st_1_1_cse
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
        & while_stage_0_3))) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01)
        & rva_in_PopNB_mioi_return_rsc_z_mxwt & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]))
        & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))
        & rva_in_reg_rw_and_5_cse ) begin
      pe_config_output_counter_sva_dfm_1 <= MUX_v_8_2_2(8'b00000000, pe_config_output_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1441_tmp ) begin
      pe_config_input_counter_sva_dfm_1 <= MUX_v_8_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl,
          PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_1_nl,
          rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_mux_27_itm_1 <= 1'b0;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= 4'b0000;
      weight_write_data_data_0_15_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_14_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_13_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_12_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_11_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_10_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_9_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_8_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= 11'b00000000000;
    end
    else if ( while_if_and_15_cse ) begin
      while_if_mux_27_itm_1 <= MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_27_nl,
          rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:0])
          & ({{3{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_4_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
      weight_write_data_data_0_15_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:120])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_14_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[119:112])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_13_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:104])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_12_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[103:96])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_11_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:88])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_10_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[87:80])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_9_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:72])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_8_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:4])
          & ({{10{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_11_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_277 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_6)
        ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_4 <= 1'b0;
      rva_in_reg_rw_sva_st_4 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_6_cse ) begin
      rva_in_reg_rw_sva_st_1_4 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1;
      rva_in_reg_rw_sva_st_4 <= rva_in_reg_rw_sva_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_7 <= 1'b0;
      rva_in_reg_rw_sva_st_7 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_7_cse ) begin
      rva_in_reg_rw_sva_st_1_7 <= rva_in_reg_rw_sva_st_1_6;
      rva_in_reg_rw_sva_st_7 <= rva_in_reg_rw_sva_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_9 <= 1'b0;
      rva_in_reg_rw_sva_st_9 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_8_cse ) begin
      rva_in_reg_rw_sva_st_1_9 <= rva_in_reg_rw_sva_st_1_8;
      rva_in_reg_rw_sva_st_9 <= rva_in_reg_rw_sva_st_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= 4'b0000;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= 1'b0;
    end
    else if ( while_if_and_16_cse ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16];
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= (pe_config_num_output_sva[7]) & (~(and_319_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1))
          & PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_398_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_401_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_135_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_142_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_55_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_132_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_405_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= MUX_v_3_2_2((weight_read_addrs_1_lpi_1_dfm_1[2:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_90 & weight_mem_run_3_for_weight_mem_run_3_for_and_1_tmp
        ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_13_itm_1
          <= ~((weight_read_addrs_1_lpi_1_dfm_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2
          <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_144_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b101)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_120_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b011)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_90_itm_1 <= (pe_manager_base_weight_sva[2])
          & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_80_itm_1 <= (pe_manager_base_weight_sva[1])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 & (~
          (pe_manager_base_weight_sva[2])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1
          <= ~((pe_manager_base_weight_sva[2:1]!=2'b00) | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1 <= (pe_manager_base_weight_sva[2])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1 & (pe_manager_base_weight_sva[0])
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1
          & (pe_manager_base_weight_sva[1:0]==2'b10) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1 <= (pe_manager_base_weight_sva[2])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 & (~
          (pe_manager_base_weight_sva[1])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_233_itm_1 & (~
          (pe_manager_base_weight_sva[1])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1
          <= ~(pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1 |
          (pe_manager_base_weight_sva[1:0]!=2'b00));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_130_itm_1
          & (pe_manager_base_weight_sva[0]) & (~ (pe_manager_base_weight_sva[2]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_146_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_115_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1,
          PECore_UpdateFSM_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1,
          PECore_RunFSM_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_95_nl & while_stage_0_5 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          input_read_req_valid_lpi_1_dfm_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1 <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd
          <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_6 <=
          1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd
          <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_1
          <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_4_3 <=
          2'b00;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_2_0 <=
          3'b000;
    end
    else if ( weight_port_read_out_data_and_174_cse ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1 <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1[0];
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd
          <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1 <= reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1[0];
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1 <= reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_2[0];
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_6 <=
          reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd
          <= reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_rsp_0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_1
          <= reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_rsp_1;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_4_3 <=
          reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_1;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_2_0 <=
          reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_2[3:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_9_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1
          <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_220_enex5 ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1
          <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1[6:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_51_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_52_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_53_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_54_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_16_0_sva_dfm_1_1 <= 17'b00000000000000000;
      act_port_reg_data_176_160_sva_dfm_1_1 <= 17'b00000000000000000;
      act_port_reg_data_208_192_sva_dfm_1_1 <= 17'b00000000000000000;
      act_port_reg_data_240_224_sva_dfm_1_1 <= 17'b00000000000000000;
    end
    else if ( and_1446_cse ) begin
      act_port_reg_data_16_0_sva_dfm_1_1 <= MUX1HOT_v_17_3_2((readslicef_28_17_11(PECore_RunScale_if_for_1_scaled_val_mul_1_nl)),
          Datapath_for_2_ProductSum_for_acc_2_1_16_0, act_port_reg_data_16_0_sva_dfm_3,
          {(~ or_dcpl_287) , PECore_RunMac_and_cse , PECore_RunMac_and_4_cse});
      act_port_reg_data_176_160_sva_dfm_1_1 <= MUX1HOT_v_17_3_2((readslicef_28_17_11(PECore_RunScale_if_for_6_scaled_val_mul_1_nl)),
          Datapath_for_2_ProductSum_for_acc_3_1_16_0, act_port_reg_data_176_160_sva_dfm_3,
          {(~ or_dcpl_287) , PECore_RunMac_and_cse , PECore_RunMac_and_4_cse});
      act_port_reg_data_208_192_sva_dfm_1_1 <= MUX1HOT_v_17_3_2((readslicef_28_17_11(PECore_RunScale_if_for_7_scaled_val_mul_1_nl)),
          Datapath_for_4_ProductSum_for_acc_2_1_16_0, act_port_reg_data_208_192_sva_dfm_3,
          {(~ or_dcpl_287) , PECore_RunMac_and_cse , PECore_RunMac_and_4_cse});
      act_port_reg_data_240_224_sva_dfm_1_1 <= MUX1HOT_v_17_3_2((readslicef_28_17_11(PECore_RunScale_if_for_8_scaled_val_mul_1_nl)),
          Datapath_for_4_ProductSum_for_acc_3_1_16_0, act_port_reg_data_240_224_sva_dfm_3,
          {(~ or_dcpl_287) , PECore_RunMac_and_cse , PECore_RunMac_and_4_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_2_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & and_dcpl_90 & weight_mem_run_3_for_weight_mem_run_3_for_and_6_tmp
        ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_9 <= 1'b0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd <= 1'b0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1 <= 3'b000;
      rva_out_reg_data_47_sva_dfm_4_4 <= 1'b0;
      rva_out_reg_data_63_sva_dfm_4_4 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_4_4_7 <= 1'b0;
      rva_out_reg_data_87_80_sva_dfm_4_4_7 <= 1'b0;
      rva_out_reg_data_119_112_sva_dfm_4_4_7 <= 1'b0;
      rva_out_reg_data_111_104_sva_dfm_4_4_7 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_4_4_6 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_4_4_5_4 <= 2'b00;
    end
    else if ( input_read_req_valid_and_1_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_9 <= input_read_req_valid_lpi_1_dfm_1_8;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd <= rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1;
      rva_out_reg_data_47_sva_dfm_4_4 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      rva_out_reg_data_63_sva_dfm_4_4 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
      rva_out_reg_data_95_88_sva_dfm_4_4_7 <= reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd;
      rva_out_reg_data_87_80_sva_dfm_4_4_7 <= reg_rva_out_reg_data_87_80_sva_dfm_4_3_ftd;
      rva_out_reg_data_119_112_sva_dfm_4_4_7 <= reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd;
      rva_out_reg_data_111_104_sva_dfm_4_4_7 <= reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd;
      rva_out_reg_data_95_88_sva_dfm_4_4_6 <= reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_0;
      rva_out_reg_data_95_88_sva_dfm_4_4_5_4 <= reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_7_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_157_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= rva_out_reg_data_30_25_sva_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_7 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_158_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_7 <= rva_out_reg_data_23_17_sva_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_159_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= rva_out_reg_data_15_9_sva_dfm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_160_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= rva_out_reg_data_35_32_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_161_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_4 <= rva_out_reg_data_46_40_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_162_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_4 <= rva_out_reg_data_62_56_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_163_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_4 <= rva_out_reg_data_55_48_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_120_sva_dfm_4_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_164_enex5 ) begin
      rva_out_reg_data_127_120_sva_dfm_4_4 <= rva_out_reg_data_127_120_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_165_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd <= rva_out_reg_data_103_96_sva_dfm_4_3_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_166_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_103_96_sva_dfm_4_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_72_sva_dfm_4_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_167_enex5 ) begin
      rva_out_reg_data_79_72_sva_dfm_4_4 <= rva_out_reg_data_79_72_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_4_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_168_enex5 ) begin
      rva_out_reg_data_71_64_sva_dfm_4_4 <= rva_out_reg_data_71_64_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Datapath_for_2_ProductSum_for_acc_2_1_17 <= 1'b0;
      Datapath_for_2_ProductSum_for_acc_3_1_17 <= 1'b0;
      Datapath_for_4_ProductSum_for_acc_2_1_17 <= 1'b0;
      Datapath_for_4_ProductSum_for_acc_3_1_17 <= 1'b0;
    end
    else if ( ProductSum_for_and_cse ) begin
      Datapath_for_2_ProductSum_for_acc_2_1_17 <= Datapath_for_4_ProductSum_for_acc_9_cmp_31_z[17];
      Datapath_for_2_ProductSum_for_acc_3_1_17 <= Datapath_for_4_ProductSum_for_acc_9_cmp_30_z[17];
      Datapath_for_4_ProductSum_for_acc_2_1_17 <= Datapath_for_4_ProductSum_for_acc_9_cmp_63_z[17];
      Datapath_for_4_ProductSum_for_acc_3_1_17 <= Datapath_for_4_ProductSum_for_acc_9_cmp_62_z[17];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Datapath_for_2_ProductSum_for_acc_2_1_16_0 <= 17'b00000000000000000;
      Datapath_for_2_ProductSum_for_acc_3_1_16_0 <= 17'b00000000000000000;
      Datapath_for_4_ProductSum_for_acc_2_1_16_0 <= 17'b00000000000000000;
      Datapath_for_4_ProductSum_for_acc_3_1_16_0 <= 17'b00000000000000000;
    end
    else if ( and_1464_cse ) begin
      Datapath_for_2_ProductSum_for_acc_2_1_16_0 <= MUX_v_17_2_2(act_port_reg_operator_for_act_port_reg_operator_for_and_nl,
          (Datapath_for_4_ProductSum_for_acc_9_cmp_31_z[16:0]), ProductSum_for_and_8_cse);
      Datapath_for_2_ProductSum_for_acc_3_1_16_0 <= MUX_v_17_2_2(act_port_reg_operator_for_act_port_reg_operator_for_and_1_nl,
          (Datapath_for_4_ProductSum_for_acc_9_cmp_30_z[16:0]), ProductSum_for_and_8_cse);
      Datapath_for_4_ProductSum_for_acc_2_1_16_0 <= MUX_v_17_2_2(act_port_reg_operator_for_act_port_reg_operator_for_and_2_nl,
          (Datapath_for_4_ProductSum_for_acc_9_cmp_63_z[16:0]), ProductSum_for_and_8_cse);
      Datapath_for_4_ProductSum_for_acc_3_1_16_0 <= MUX_v_17_2_2(act_port_reg_operator_for_act_port_reg_operator_for_and_3_nl,
          (Datapath_for_4_ProductSum_for_acc_9_cmp_62_z[16:0]), ProductSum_for_and_8_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_acc_40_itm_1 <= 20'b00000000000000000000;
      ProductSum_for_acc_41_itm_1 <= 19'b0000000000000000000;
      ProductSum_for_acc_24_itm_1 <= 20'b00000000000000000000;
      ProductSum_for_acc_25_itm_1 <= 19'b0000000000000000000;
    end
    else if ( ProductSum_for_and_2_cse ) begin
      ProductSum_for_acc_40_itm_1 <= nl_ProductSum_for_acc_40_itm_1[19:0];
      ProductSum_for_acc_41_itm_1 <= nl_ProductSum_for_acc_41_itm_1[18:0];
      ProductSum_for_acc_24_itm_1 <= nl_ProductSum_for_acc_24_itm_1[19:0];
      ProductSum_for_acc_25_itm_1 <= nl_ProductSum_for_acc_25_itm_1[18:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd <= 1'b0;
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_1 <= 2'b00;
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= 1'b0;
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_rsp_0 <= 1'b0;
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_rsp_1 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_182_ssc ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd <= weight_port_read_out_data_0_1_sva_dfm_2_rsp_0;
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_1 <= weight_port_read_out_data_0_2_sva_dfm_2_rsp_1;
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_0_sva_dfm_2_7;
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_rsp_0 <= weight_port_read_out_data_0_2_sva_dfm_2_rsp_0_1;
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_rsp_1 <= weight_port_read_out_data_0_2_sva_dfm_2_rsp_0_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_221_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1 <= weight_port_read_out_data_0_1_sva_dfm_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_2 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_222_enex5 ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_ftd_2 <= weight_port_read_out_data_0_2_sva_dfm_2_rsp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_19_0_sva <= 20'b00000000000000000000;
      accum_vector_data_0_19_0_sva <= 20'b00000000000000000000;
      accum_vector_data_6_19_0_sva <= 20'b00000000000000000000;
      accum_vector_data_5_19_0_sva <= 20'b00000000000000000000;
    end
    else if ( and_1476_cse ) begin
      accum_vector_data_7_19_0_sva <= MUX_v_20_2_2(20'b00000000000000000000, ProductSum_for_acc_nl,
          PECore_UpdateFSM_switch_lp_not_37_nl);
      accum_vector_data_0_19_0_sva <= MUX_v_20_2_2(20'b00000000000000000000, ProductSum_for_acc_46_nl,
          PECore_UpdateFSM_switch_lp_not_23_nl);
      accum_vector_data_6_19_0_sva <= MUX_v_20_2_2(20'b00000000000000000000, ProductSum_for_acc_42_nl,
          PECore_UpdateFSM_switch_lp_not_38_nl);
      accum_vector_data_5_19_0_sva <= MUX_v_20_2_2(20'b00000000000000000000, ProductSum_for_acc_34_nl,
          PECore_UpdateFSM_switch_lp_not_39_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_3_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= 8'b00000000;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_empty_and_enex5 ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= weight_mem_write_arbxbar_xbar_for_empty_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_data_sva_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rva_in_reg_data_and_tmp ) begin
      rva_in_reg_data_sva_1 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_33 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_5)
        ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_6 <= 1'b0;
      rva_in_reg_rw_sva_st_6 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_11_cse ) begin
      rva_in_reg_rw_sva_st_1_6 <= rva_in_reg_rw_sva_st_1_5;
      rva_in_reg_rw_sva_st_6 <= rva_in_reg_rw_sva_st_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_1 <= 2'b00;
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= 1'b0;
    end
    else if ( pe_manager_base_weight_and_6_cse ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_1 <= pe_manager_base_weight_sva[1:0];
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= weight_read_addrs_4_14_2_lpi_1_dfm_1[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_1 <= 1'b0;
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( pe_manager_base_weight_and_7_cse ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_1 <= pe_manager_base_weight_sva[0];
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_18_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_55_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_56_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_57_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_58_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= 1'b0;
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd <= 1'b0;
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd <= 1'b0;
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd <= 1'b0;
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_ftd <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1 <= 3'b000;
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_0 <= 1'b0;
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_1 <= 2'b00;
    end
    else if ( input_read_req_valid_and_2_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= input_read_req_valid_lpi_1_dfm_1_7;
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd <= rva_out_reg_data_119_112_sva_dfm_4_2_rsp_0;
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd <= rva_out_reg_data_111_104_sva_dfm_4_2_rsp_0;
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd <= rva_out_reg_data_95_88_sva_dfm_4_2_rsp_0;
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_ftd <= rva_out_reg_data_87_80_sva_dfm_4_2_rsp_0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_39_36_sva_dfm_4_2_3;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_39_36_sva_dfm_4_2_2_0;
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_0 <= rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_6;
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_1 <= rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_5_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_11_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_6 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_169_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_6 <= rva_out_reg_data_30_25_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_6 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_170_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_6 <= rva_out_reg_data_23_17_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_171_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= rva_out_reg_data_15_9_sva_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_223_enex5 ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd <= weight_port_read_out_data_0_3_sva_dfm_2_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_224_enex5 ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd_1 <= weight_port_read_out_data_0_3_sva_dfm_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_172_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= rva_out_reg_data_35_32_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_173_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3 <= rva_out_reg_data_46_40_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_174_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_3 <= rva_out_reg_data_62_56_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_175_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3 <= rva_out_reg_data_55_48_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_120_sva_dfm_4_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_176_enex5 ) begin
      rva_out_reg_data_127_120_sva_dfm_4_3 <= rva_out_reg_data_127_120_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_177_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd_1 <= rva_out_reg_data_119_112_sva_dfm_4_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_178_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd_1 <= rva_out_reg_data_111_104_sva_dfm_4_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_ftd_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_179_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_ftd_1 <= rva_out_reg_data_87_80_sva_dfm_4_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_72_sva_dfm_4_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_180_enex5 ) begin
      rva_out_reg_data_79_72_sva_dfm_4_3 <= rva_out_reg_data_79_72_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_4_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_181_enex5 ) begin
      rva_out_reg_data_71_64_sva_dfm_4_3 <= rva_out_reg_data_71_64_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
        & while_stage_0_6 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_6_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_27_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_59_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_60_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= weight_port_read_out_data_0_0_sva_dfm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_61_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_62_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= MUX_v_128_256_2(input_mem_banks_bank_a_0_sva_dfm_2,
          input_mem_banks_bank_a_1_sva_dfm_2, input_mem_banks_bank_a_2_sva_dfm_2,
          input_mem_banks_bank_a_3_sva_dfm_2, input_mem_banks_bank_a_4_sva_dfm_2,
          input_mem_banks_bank_a_5_sva_dfm_2, input_mem_banks_bank_a_6_sva_dfm_2,
          input_mem_banks_bank_a_7_sva_dfm_2, input_mem_banks_bank_a_8_sva_dfm_2,
          input_mem_banks_bank_a_9_sva_dfm_2, input_mem_banks_bank_a_10_sva_dfm_2,
          input_mem_banks_bank_a_11_sva_dfm_2, input_mem_banks_bank_a_12_sva_dfm_2,
          input_mem_banks_bank_a_13_sva_dfm_2, input_mem_banks_bank_a_14_sva_dfm_2,
          input_mem_banks_bank_a_15_sva_dfm_2, input_mem_banks_bank_a_16_sva_dfm_2,
          input_mem_banks_bank_a_17_sva_dfm_2, input_mem_banks_bank_a_18_sva_dfm_2,
          input_mem_banks_bank_a_19_sva_dfm_2, input_mem_banks_bank_a_20_sva_dfm_2,
          input_mem_banks_bank_a_21_sva_dfm_2, input_mem_banks_bank_a_22_sva_dfm_2,
          input_mem_banks_bank_a_23_sva_dfm_2, input_mem_banks_bank_a_24_sva_dfm_2,
          input_mem_banks_bank_a_25_sva_dfm_2, input_mem_banks_bank_a_26_sva_dfm_2,
          input_mem_banks_bank_a_27_sva_dfm_2, input_mem_banks_bank_a_28_sva_dfm_2,
          input_mem_banks_bank_a_29_sva_dfm_2, input_mem_banks_bank_a_30_sva_dfm_2,
          input_mem_banks_bank_a_31_sva_dfm_2, input_mem_banks_bank_a_32_sva_dfm_2,
          input_mem_banks_bank_a_33_sva_dfm_2, input_mem_banks_bank_a_34_sva_dfm_2,
          input_mem_banks_bank_a_35_sva_dfm_2, input_mem_banks_bank_a_36_sva_dfm_2,
          input_mem_banks_bank_a_37_sva_dfm_2, input_mem_banks_bank_a_38_sva_dfm_2,
          input_mem_banks_bank_a_39_sva_dfm_2, input_mem_banks_bank_a_40_sva_dfm_2,
          input_mem_banks_bank_a_41_sva_dfm_2, input_mem_banks_bank_a_42_sva_dfm_2,
          input_mem_banks_bank_a_43_sva_dfm_2, input_mem_banks_bank_a_44_sva_dfm_2,
          input_mem_banks_bank_a_45_sva_dfm_2, input_mem_banks_bank_a_46_sva_dfm_2,
          input_mem_banks_bank_a_47_sva_dfm_2, input_mem_banks_bank_a_48_sva_dfm_2,
          input_mem_banks_bank_a_49_sva_dfm_2, input_mem_banks_bank_a_50_sva_dfm_2,
          input_mem_banks_bank_a_51_sva_dfm_2, input_mem_banks_bank_a_52_sva_dfm_2,
          input_mem_banks_bank_a_53_sva_dfm_2, input_mem_banks_bank_a_54_sva_dfm_2,
          input_mem_banks_bank_a_55_sva_dfm_2, input_mem_banks_bank_a_56_sva_dfm_2,
          input_mem_banks_bank_a_57_sva_dfm_2, input_mem_banks_bank_a_58_sva_dfm_2,
          input_mem_banks_bank_a_59_sva_dfm_2, input_mem_banks_bank_a_60_sva_dfm_2,
          input_mem_banks_bank_a_61_sva_dfm_2, input_mem_banks_bank_a_62_sva_dfm_2,
          input_mem_banks_bank_a_63_sva_dfm_2, input_mem_banks_bank_a_64_sva_dfm_2,
          input_mem_banks_bank_a_65_sva_dfm_2, input_mem_banks_bank_a_66_sva_dfm_2,
          input_mem_banks_bank_a_67_sva_dfm_2, input_mem_banks_bank_a_68_sva_dfm_2,
          input_mem_banks_bank_a_69_sva_dfm_2, input_mem_banks_bank_a_70_sva_dfm_2,
          input_mem_banks_bank_a_71_sva_dfm_2, input_mem_banks_bank_a_72_sva_dfm_2,
          input_mem_banks_bank_a_73_sva_dfm_2, input_mem_banks_bank_a_74_sva_dfm_2,
          input_mem_banks_bank_a_75_sva_dfm_2, input_mem_banks_bank_a_76_sva_dfm_2,
          input_mem_banks_bank_a_77_sva_dfm_2, input_mem_banks_bank_a_78_sva_dfm_2,
          input_mem_banks_bank_a_79_sva_dfm_2, input_mem_banks_bank_a_80_sva_dfm_2,
          input_mem_banks_bank_a_81_sva_dfm_2, input_mem_banks_bank_a_82_sva_dfm_2,
          input_mem_banks_bank_a_83_sva_dfm_2, input_mem_banks_bank_a_84_sva_dfm_2,
          input_mem_banks_bank_a_85_sva_dfm_2, input_mem_banks_bank_a_86_sva_dfm_2,
          input_mem_banks_bank_a_87_sva_dfm_2, input_mem_banks_bank_a_88_sva_dfm_2,
          input_mem_banks_bank_a_89_sva_dfm_2, input_mem_banks_bank_a_90_sva_dfm_2,
          input_mem_banks_bank_a_91_sva_dfm_2, input_mem_banks_bank_a_92_sva_dfm_2,
          input_mem_banks_bank_a_93_sva_dfm_2, input_mem_banks_bank_a_94_sva_dfm_2,
          input_mem_banks_bank_a_95_sva_dfm_2, input_mem_banks_bank_a_96_sva_dfm_2,
          input_mem_banks_bank_a_97_sva_dfm_2, input_mem_banks_bank_a_98_sva_dfm_2,
          input_mem_banks_bank_a_99_sva_dfm_2, input_mem_banks_bank_a_100_sva_dfm_2,
          input_mem_banks_bank_a_101_sva_dfm_2, input_mem_banks_bank_a_102_sva_dfm_2,
          input_mem_banks_bank_a_103_sva_dfm_2, input_mem_banks_bank_a_104_sva_dfm_2,
          input_mem_banks_bank_a_105_sva_dfm_2, input_mem_banks_bank_a_106_sva_dfm_2,
          input_mem_banks_bank_a_107_sva_dfm_2, input_mem_banks_bank_a_108_sva_dfm_2,
          input_mem_banks_bank_a_109_sva_dfm_2, input_mem_banks_bank_a_110_sva_dfm_2,
          input_mem_banks_bank_a_111_sva_dfm_2, input_mem_banks_bank_a_112_sva_dfm_2,
          input_mem_banks_bank_a_113_sva_dfm_2, input_mem_banks_bank_a_114_sva_dfm_2,
          input_mem_banks_bank_a_115_sva_dfm_2, input_mem_banks_bank_a_116_sva_dfm_2,
          input_mem_banks_bank_a_117_sva_dfm_2, input_mem_banks_bank_a_118_sva_dfm_2,
          input_mem_banks_bank_a_119_sva_dfm_2, input_mem_banks_bank_a_120_sva_dfm_2,
          input_mem_banks_bank_a_121_sva_dfm_2, input_mem_banks_bank_a_122_sva_dfm_2,
          input_mem_banks_bank_a_123_sva_dfm_2, input_mem_banks_bank_a_124_sva_dfm_2,
          input_mem_banks_bank_a_125_sva_dfm_2, input_mem_banks_bank_a_126_sva_dfm_2,
          input_mem_banks_bank_a_127_sva_dfm_2, input_mem_banks_bank_a_128_sva_dfm_2,
          input_mem_banks_bank_a_129_sva_dfm_2, input_mem_banks_bank_a_130_sva_dfm_2,
          input_mem_banks_bank_a_131_sva_dfm_2, input_mem_banks_bank_a_132_sva_dfm_2,
          input_mem_banks_bank_a_133_sva_dfm_2, input_mem_banks_bank_a_134_sva_dfm_2,
          input_mem_banks_bank_a_135_sva_dfm_2, input_mem_banks_bank_a_136_sva_dfm_2,
          input_mem_banks_bank_a_137_sva_dfm_2, input_mem_banks_bank_a_138_sva_dfm_2,
          input_mem_banks_bank_a_139_sva_dfm_2, input_mem_banks_bank_a_140_sva_dfm_2,
          input_mem_banks_bank_a_141_sva_dfm_2, input_mem_banks_bank_a_142_sva_dfm_2,
          input_mem_banks_bank_a_143_sva_dfm_2, input_mem_banks_bank_a_144_sva_dfm_2,
          input_mem_banks_bank_a_145_sva_dfm_2, input_mem_banks_bank_a_146_sva_dfm_2,
          input_mem_banks_bank_a_147_sva_dfm_2, input_mem_banks_bank_a_148_sva_dfm_2,
          input_mem_banks_bank_a_149_sva_dfm_2, input_mem_banks_bank_a_150_sva_dfm_2,
          input_mem_banks_bank_a_151_sva_dfm_2, input_mem_banks_bank_a_152_sva_dfm_2,
          input_mem_banks_bank_a_153_sva_dfm_2, input_mem_banks_bank_a_154_sva_dfm_2,
          input_mem_banks_bank_a_155_sva_dfm_2, input_mem_banks_bank_a_156_sva_dfm_2,
          input_mem_banks_bank_a_157_sva_dfm_2, input_mem_banks_bank_a_158_sva_dfm_2,
          input_mem_banks_bank_a_159_sva_dfm_2, input_mem_banks_bank_a_160_sva_dfm_2,
          input_mem_banks_bank_a_161_sva_dfm_2, input_mem_banks_bank_a_162_sva_dfm_2,
          input_mem_banks_bank_a_163_sva_dfm_2, input_mem_banks_bank_a_164_sva_dfm_2,
          input_mem_banks_bank_a_165_sva_dfm_2, input_mem_banks_bank_a_166_sva_dfm_2,
          input_mem_banks_bank_a_167_sva_dfm_2, input_mem_banks_bank_a_168_sva_dfm_2,
          input_mem_banks_bank_a_169_sva_dfm_2, input_mem_banks_bank_a_170_sva_dfm_2,
          input_mem_banks_bank_a_171_sva_dfm_2, input_mem_banks_bank_a_172_sva_dfm_2,
          input_mem_banks_bank_a_173_sva_dfm_2, input_mem_banks_bank_a_174_sva_dfm_2,
          input_mem_banks_bank_a_175_sva_dfm_2, input_mem_banks_bank_a_176_sva_dfm_2,
          input_mem_banks_bank_a_177_sva_dfm_2, input_mem_banks_bank_a_178_sva_dfm_2,
          input_mem_banks_bank_a_179_sva_dfm_2, input_mem_banks_bank_a_180_sva_dfm_2,
          input_mem_banks_bank_a_181_sva_dfm_2, input_mem_banks_bank_a_182_sva_dfm_2,
          input_mem_banks_bank_a_183_sva_dfm_2, input_mem_banks_bank_a_184_sva_dfm_2,
          input_mem_banks_bank_a_185_sva_dfm_2, input_mem_banks_bank_a_186_sva_dfm_2,
          input_mem_banks_bank_a_187_sva_dfm_2, input_mem_banks_bank_a_188_sva_dfm_2,
          input_mem_banks_bank_a_189_sva_dfm_2, input_mem_banks_bank_a_190_sva_dfm_2,
          input_mem_banks_bank_a_191_sva_dfm_2, input_mem_banks_bank_a_192_sva_dfm_2,
          input_mem_banks_bank_a_193_sva_dfm_2, input_mem_banks_bank_a_194_sva_dfm_2,
          input_mem_banks_bank_a_195_sva_dfm_2, input_mem_banks_bank_a_196_sva_dfm_2,
          input_mem_banks_bank_a_197_sva_dfm_2, input_mem_banks_bank_a_198_sva_dfm_2,
          input_mem_banks_bank_a_199_sva_dfm_2, input_mem_banks_bank_a_200_sva_dfm_2,
          input_mem_banks_bank_a_201_sva_dfm_2, input_mem_banks_bank_a_202_sva_dfm_2,
          input_mem_banks_bank_a_203_sva_dfm_2, input_mem_banks_bank_a_204_sva_dfm_2,
          input_mem_banks_bank_a_205_sva_dfm_2, input_mem_banks_bank_a_206_sva_dfm_2,
          input_mem_banks_bank_a_207_sva_dfm_2, input_mem_banks_bank_a_208_sva_dfm_2,
          input_mem_banks_bank_a_209_sva_dfm_2, input_mem_banks_bank_a_210_sva_dfm_2,
          input_mem_banks_bank_a_211_sva_dfm_2, input_mem_banks_bank_a_212_sva_dfm_2,
          input_mem_banks_bank_a_213_sva_dfm_2, input_mem_banks_bank_a_214_sva_dfm_2,
          input_mem_banks_bank_a_215_sva_dfm_2, input_mem_banks_bank_a_216_sva_dfm_2,
          input_mem_banks_bank_a_217_sva_dfm_2, input_mem_banks_bank_a_218_sva_dfm_2,
          input_mem_banks_bank_a_219_sva_dfm_2, input_mem_banks_bank_a_220_sva_dfm_2,
          input_mem_banks_bank_a_221_sva_dfm_2, input_mem_banks_bank_a_222_sva_dfm_2,
          input_mem_banks_bank_a_223_sva_dfm_2, input_mem_banks_bank_a_224_sva_dfm_2,
          input_mem_banks_bank_a_225_sva_dfm_2, input_mem_banks_bank_a_226_sva_dfm_2,
          input_mem_banks_bank_a_227_sva_dfm_2, input_mem_banks_bank_a_228_sva_dfm_2,
          input_mem_banks_bank_a_229_sva_dfm_2, input_mem_banks_bank_a_230_sva_dfm_2,
          input_mem_banks_bank_a_231_sva_dfm_2, input_mem_banks_bank_a_232_sva_dfm_2,
          input_mem_banks_bank_a_233_sva_dfm_2, input_mem_banks_bank_a_234_sva_dfm_2,
          input_mem_banks_bank_a_235_sva_dfm_2, input_mem_banks_bank_a_236_sva_dfm_2,
          input_mem_banks_bank_a_237_sva_dfm_2, input_mem_banks_bank_a_238_sva_dfm_2,
          input_mem_banks_bank_a_239_sva_dfm_2, input_mem_banks_bank_a_240_sva_dfm_2,
          input_mem_banks_bank_a_241_sva_dfm_2, input_mem_banks_bank_a_242_sva_dfm_2,
          input_mem_banks_bank_a_243_sva_dfm_2, input_mem_banks_bank_a_244_sva_dfm_2,
          input_mem_banks_bank_a_245_sva_dfm_2, input_mem_banks_bank_a_246_sva_dfm_2,
          input_mem_banks_bank_a_247_sva_dfm_2, input_mem_banks_bank_a_248_sva_dfm_2,
          input_mem_banks_bank_a_249_sva_dfm_2, input_mem_banks_bank_a_250_sva_dfm_2,
          input_mem_banks_bank_a_251_sva_dfm_2, input_mem_banks_bank_a_252_sva_dfm_2,
          input_mem_banks_bank_a_253_sva_dfm_2, input_mem_banks_bank_a_254_sva_dfm_2,
          input_mem_banks_bank_a_255_sva_dfm_2, input_mem_banks_read_1_for_mux_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_2_3 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_2_2_0 <= 3'b000;
      rva_out_reg_data_95_88_sva_dfm_4_2_rsp_0 <= 1'b0;
      rva_out_reg_data_87_80_sva_dfm_4_2_rsp_0 <= 1'b0;
      rva_out_reg_data_119_112_sva_dfm_4_2_rsp_0 <= 1'b0;
      rva_out_reg_data_111_104_sva_dfm_4_2_rsp_0 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_6 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_5_4 <= 2'b00;
    end
    else if ( input_read_req_valid_and_3_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= input_read_req_valid_lpi_1_dfm_1_6;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
      rva_out_reg_data_39_36_sva_dfm_4_2_3 <= rva_out_reg_data_39_36_sva_dfm_4_1_3;
      rva_out_reg_data_39_36_sva_dfm_4_2_2_0 <= rva_out_reg_data_39_36_sva_dfm_4_1_2_0;
      rva_out_reg_data_95_88_sva_dfm_4_2_rsp_0 <= rva_out_reg_data_95_88_sva_dfm_4_1_7;
      rva_out_reg_data_87_80_sva_dfm_4_2_rsp_0 <= rva_out_reg_data_87_80_sva_dfm_4_1_7;
      rva_out_reg_data_119_112_sva_dfm_4_2_rsp_0 <= rva_out_reg_data_119_112_sva_dfm_4_1_7;
      rva_out_reg_data_111_104_sva_dfm_4_2_rsp_0 <= rva_out_reg_data_111_104_sva_dfm_4_1_7;
      rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_6 <= reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd;
      rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_5_4 <= reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_15_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_182_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= rva_out_reg_data_30_25_sva_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_183_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= rva_out_reg_data_23_17_sva_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_7 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_184_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_7 <= rva_out_reg_data_15_9_sva_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_185_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= rva_out_reg_data_35_32_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_186_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2 <= rva_out_reg_data_46_40_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_187_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_2 <= rva_out_reg_data_62_56_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_188_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2 <= rva_out_reg_data_55_48_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_120_sva_dfm_4_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_189_enex5 ) begin
      rva_out_reg_data_127_120_sva_dfm_4_2 <= rva_out_reg_data_127_120_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_72_sva_dfm_4_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_190_enex5 ) begin
      rva_out_reg_data_79_72_sva_dfm_4_2 <= rva_out_reg_data_79_72_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_4_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_191_enex5 ) begin
      rva_out_reg_data_71_64_sva_dfm_4_2 <= rva_out_reg_data_71_64_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_6_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_221_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_221_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_225_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_225_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_229_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_229_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_233_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_233_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_237_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_237_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_241_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_241_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_245_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_245_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_249_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_249_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_253_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_253_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_257_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_257_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_261_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_261_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_265_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_265_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_269_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_269_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_273_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_273_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_277_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_277_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_281_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_281_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_285_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_285_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_289_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_289_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_293_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_293_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_297_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_297_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_301_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_301_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_305_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_305_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_309_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_309_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_313_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_313_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_317_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_317_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_321_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_321_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_325_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_325_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_329_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_329_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_333_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_333_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_337_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_337_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_341_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_341_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_345_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_345_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_349_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_349_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_353_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_353_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_357_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_357_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_361_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_361_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_365_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_365_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_369_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_369_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_373_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_373_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_377_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_377_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_381_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_381_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_385_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_385_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_389_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_389_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_393_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_393_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_397_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_397_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_401_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_401_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_405_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_405_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_409_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_409_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_413_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_413_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_417_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_417_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_421_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_421_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_425_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_425_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_429_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_429_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_433_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_433_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_437_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_437_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_441_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_441_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_445_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_445_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_449_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_449_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_453_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_453_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_457_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_457_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_461_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_461_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_465_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_465_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_469_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_469_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_473_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_473_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_477_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_477_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_481_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_481_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_485_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_485_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_489_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_489_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_493_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_493_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_497_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_497_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_501_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_501_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_505_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_505_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_509_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_509_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_513_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_513_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_517_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_517_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_521_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_521_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_525_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_525_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_529_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_529_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_533_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_533_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_537_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_537_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_541_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_541_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_545_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_545_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_549_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_549_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_553_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_553_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_557_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_557_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_561_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_561_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_565_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_565_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_569_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_569_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_573_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_573_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_577_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_577_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_581_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_581_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_585_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_585_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_589_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_589_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_593_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_593_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_597_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_597_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_601_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_601_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_605_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_605_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_609_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_609_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_613_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_613_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_617_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_617_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_621_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_621_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_625_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_625_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_629_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_629_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_633_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_633_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_637_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_637_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_641_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_641_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_645_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_645_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_649_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_649_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_653_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_653_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_657_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_657_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_661_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_661_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_665_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_665_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_669_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_669_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_673_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_673_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_677_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_677_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_681_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_681_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_685_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_685_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_689_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_689_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_693_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_693_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_697_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_697_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_701_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_701_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_705_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_705_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_709_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_709_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_713_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_713_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_717_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_717_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_721_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_721_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_725_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_725_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_729_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_729_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_733_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_733_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_737_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_737_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_741_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_741_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_745_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_745_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_749_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_749_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_753_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_753_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_757_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_757_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_761_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_761_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_765_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_765_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_769_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_769_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_773_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_773_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_777_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_777_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_781_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_781_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_785_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_785_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_789_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_789_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_793_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_793_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_797_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_797_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_801_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_801_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_805_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_805_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_809_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_809_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_813_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_813_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_817_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_817_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_821_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_821_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_825_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_825_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_829_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_829_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_833_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_833_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_837_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_837_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_841_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_841_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_845_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_845_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_849_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_849_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_853_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_853_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_857_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_857_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_861_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_861_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_865_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_865_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_869_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_869_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_873_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_873_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_877_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_877_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_881_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_881_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_885_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_885_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_889_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_889_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_893_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_893_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_897_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_897_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_901_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_901_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_905_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_905_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_909_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_909_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_913_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_913_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_917_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_917_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_921_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_921_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_925_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_925_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_929_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_929_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_933_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_933_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_937_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_937_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_941_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_941_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_945_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_945_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_949_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_949_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_953_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_953_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_957_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_957_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_961_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_961_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_965_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_965_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_969_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_969_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_973_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_973_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_977_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_977_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_981_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_981_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_985_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_985_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_989_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_989_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_993_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_993_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_997_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_997_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1001_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1001_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1005_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1005_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1009_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1009_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1013_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1013_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1017_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1017_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1021_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1021_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1025_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1025_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1029_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1029_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1033_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1033_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1037_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1037_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1041_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1041_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1045_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1045_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1049_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1049_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1053_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1053_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1057_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1057_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1061_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1061_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1065_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1065_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1069_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1069_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1073_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1073_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1077_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1077_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1081_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1081_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1085_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1085_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1089_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1089_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1093_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1093_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1097_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1097_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1101_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1101_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1105_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1105_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1109_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1109_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1113_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1113_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1117_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1117_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1121_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1121_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1125_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1125_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1129_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1129_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1133_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1133_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1137_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1137_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1141_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1141_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1145_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1145_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1149_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1149_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1153_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1153_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1157_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1157_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1161_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1161_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1165_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1165_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1169_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1169_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1173_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1173_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1177_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1177_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1181_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1181_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1185_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1185_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1189_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1189_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1193_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1193_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1197_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1197_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1201_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1201_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1205_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1205_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1209_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1209_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1213_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1213_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1217_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1217_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1221_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1221_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1225_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1225_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1229_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1229_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1233_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1233_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1237_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1237_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1241_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1241_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_36_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_4[0];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_4[8];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[16];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[31];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_63_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_64_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:17];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_65_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[30:25];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= 1'b0;
      rva_out_reg_data_79_72_sva_dfm_4_1 <= 8'b00000000;
      rva_out_reg_data_71_64_sva_dfm_4_1 <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_4_1_7 <= 1'b0;
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd <= 1'b0;
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd_1 <= 2'b00;
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd_2 <= 4'b0000;
      rva_out_reg_data_87_80_sva_dfm_4_1_7 <= 1'b0;
      rva_out_reg_data_87_80_sva_dfm_4_1_6_0 <= 7'b0000000;
    end
    else if ( input_read_req_valid_and_4_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_295_itm_1;
      rva_out_reg_data_79_72_sva_dfm_4_1 <= rva_out_reg_data_79_72_sva_dfm_7;
      rva_out_reg_data_71_64_sva_dfm_4_1 <= rva_out_reg_data_71_64_sva_dfm_7;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
      rva_out_reg_data_95_88_sva_dfm_4_1_7 <= rva_out_reg_data_95_88_sva_dfm_7_7;
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd <= rva_out_reg_data_95_88_sva_dfm_7_6;
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd_1 <= rva_out_reg_data_95_88_sva_dfm_7_5_4;
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd_2 <= rva_out_reg_data_95_88_sva_dfm_7_3_0;
      rva_out_reg_data_87_80_sva_dfm_4_1_7 <= rva_out_reg_data_87_80_sva_dfm_7_7;
      rva_out_reg_data_87_80_sva_dfm_4_1_6_0 <= rva_out_reg_data_87_80_sva_dfm_7_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_19_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_4 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_192_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_4 <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_193_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_4 <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_6 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_194_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_6 <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_4_1 <= 7'b0000000;
      rva_out_reg_data_62_56_sva_dfm_4_1 <= 7'b0000000;
      rva_out_reg_data_55_48_sva_dfm_4_1 <= 8'b00000000;
    end
    else if ( and_1489_cse ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= MUX1HOT_v_4_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_3_0,
          rva_out_reg_data_35_32_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[35:32]),
          (weight_port_read_out_data_0_4_sva_dfm_mx0w2_6_0[3:0]), {PECore_PushAxiRsp_if_asn_89
          , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_46_40_sva_dfm_4_1 <= MUX1HOT_v_7_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1_6_0,
          rva_out_reg_data_46_40_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[46:40]),
          weight_port_read_out_data_0_5_sva_dfm_mx0w2_6_0, {PECore_PushAxiRsp_if_asn_89
          , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_62_56_sva_dfm_4_1 <= MUX1HOT_v_7_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1_6_0,
          rva_out_reg_data_62_56_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[62:56]),
          (weight_port_read_out_data_0_7_sva_dfm_mx0w2[6:0]), {PECore_PushAxiRsp_if_asn_89
          , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_55_48_sva_dfm_4_1 <= MUX1HOT_v_8_4_2(rva_out_reg_data_55_48_sva_dfm_1_5,
          rva_out_reg_data_55_48_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_8_7_0_sdt_47_40_sva_1,
          {PECore_PushAxiRsp_if_asn_89 , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87
          , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_120_sva_dfm_4_1 <= 8'b00000000;
      rva_out_reg_data_119_112_sva_dfm_4_1_7 <= 1'b0;
      rva_out_reg_data_119_112_sva_dfm_4_1_6_0 <= 7'b0000000;
      rva_out_reg_data_111_104_sva_dfm_4_1_7 <= 1'b0;
      rva_out_reg_data_111_104_sva_dfm_4_1_6_0 <= 7'b0000000;
      rva_out_reg_data_103_96_sva_dfm_4_1_7_4 <= 4'b0000;
      rva_out_reg_data_103_96_sva_dfm_4_1_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_98_cse ) begin
      rva_out_reg_data_127_120_sva_dfm_4_1 <= MUX1HOT_v_8_3_2(rva_out_reg_data_127_120_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000,
          weight_port_read_out_data_4_15_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_693_nl , nor_612_nl});
      rva_out_reg_data_119_112_sva_dfm_4_1_7 <= MUX1HOT_s_1_3_2(rva_out_reg_data_119_112_sva_dfm_4_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014[7]),
          (weight_port_read_out_data_3_14_sva_dfm_1[7]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_695_ssc , nor_613_ssc});
      rva_out_reg_data_119_112_sva_dfm_4_1_6_0 <= MUX1HOT_v_7_3_2(rva_out_reg_data_119_112_sva_dfm_4_mx0w0_6_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014[6:0]),
          (weight_port_read_out_data_3_14_sva_dfm_1[6:0]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_695_ssc , nor_613_ssc});
      rva_out_reg_data_111_104_sva_dfm_4_1_7 <= MUX1HOT_s_1_3_2(rva_out_reg_data_111_104_sva_dfm_4_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000[7]),
          (weight_port_read_out_data_2_15_sva_dfm_1[7]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_697_ssc , nor_614_ssc});
      rva_out_reg_data_111_104_sva_dfm_4_1_6_0 <= MUX1HOT_v_7_3_2(rva_out_reg_data_111_104_sva_dfm_4_mx0w0_6_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_p000000[6:0]),
          (weight_port_read_out_data_2_15_sva_dfm_1[6:0]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_697_ssc , nor_614_ssc});
      rva_out_reg_data_103_96_sva_dfm_4_1_7_4 <= MUX1HOT_v_4_3_2(rva_out_reg_data_103_96_sva_dfm_4_mx0w0_7_4,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014[7:4]),
          (weight_port_read_out_data_1_14_sva_dfm_1[7:4]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_699_ssc , nor_615_ssc});
      rva_out_reg_data_103_96_sva_dfm_4_1_3_0 <= MUX1HOT_v_4_3_2(rva_out_reg_data_103_96_sva_dfm_4_mx0w0_3_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000014[3:0]),
          (weight_port_read_out_data_1_14_sva_dfm_1[3:0]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_699_ssc , nor_615_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_7_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_62_56_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_46_40_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_35_32_sva_dfm_6 <= 4'b0000;
    end
    else if ( and_1506_cse ) begin
      rva_out_reg_data_55_48_sva_dfm_6 <= rva_out_reg_data_55_48_sva_dfm_6_mx1;
      rva_out_reg_data_62_56_sva_dfm_6 <= rva_out_reg_data_62_56_sva_dfm_6_mx1;
      rva_out_reg_data_46_40_sva_dfm_6 <= rva_out_reg_data_46_40_sva_dfm_6_mx1;
      rva_out_reg_data_35_32_sva_dfm_6 <= rva_out_reg_data_35_32_sva_dfm_6_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_23_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & ((and_dcpl_41 & rva_in_reg_rw_sva_5) | PECore_PushAxiRsp_mux_23_itm_1_mx0c1)
        ) begin
      PECore_PushAxiRsp_mux_23_itm_1 <= MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
          weight_port_read_out_data_mux_144_nl, PECore_PushAxiRsp_mux_23_itm_1_mx0c1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(nand_40_cse | rva_in_reg_rw_sva_5 | (~ fsm_output)))
        ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          weight_port_read_out_data_0_5_sva_dfm_mx0w2_7, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_44_tmp ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= MUX1HOT_v_128_3_2(input_mem_banks_read_read_data_lpi_1_dfm_1_3,
          weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d, weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1,
          {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          , and_703_nl , nor_616_nl});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_5 <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7_4
          <= 4'b0000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_3_0
          <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_111_cse ) begin
      rva_out_reg_data_55_48_sva_dfm_1_5 <= MUX_v_8_2_2(rva_out_reg_data_55_48_sva_dfm_1_4,
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7_4
          <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm[7:4];
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_3_0
          <= MUX_v_4_2_2(rva_out_reg_data_39_36_sva_dfm_1_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm[3:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_79_72_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_127_120_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_87_80_sva_dfm_6_6_0 <= 7'b0000000;
      rva_out_reg_data_103_96_sva_dfm_6_7_4 <= 4'b0000;
      rva_out_reg_data_103_96_sva_dfm_6_3_0 <= 4'b0000;
      rva_out_reg_data_111_104_sva_dfm_6_6_0 <= 7'b0000000;
      rva_out_reg_data_119_112_sva_dfm_6_6_0 <= 7'b0000000;
      rva_out_reg_data_95_88_sva_dfm_6_3_0 <= 4'b0000;
    end
    else if ( and_1526_cse ) begin
      rva_out_reg_data_71_64_sva_dfm_6 <= rva_out_reg_data_71_64_sva_dfm_7;
      rva_out_reg_data_79_72_sva_dfm_6 <= rva_out_reg_data_79_72_sva_dfm_7;
      rva_out_reg_data_127_120_sva_dfm_6 <= rva_out_reg_data_127_120_sva_dfm_4_mx0w0;
      rva_out_reg_data_87_80_sva_dfm_6_6_0 <= rva_out_reg_data_87_80_sva_dfm_7_6_0;
      rva_out_reg_data_103_96_sva_dfm_6_7_4 <= rva_out_reg_data_103_96_sva_dfm_4_mx0w0_7_4;
      rva_out_reg_data_103_96_sva_dfm_6_3_0 <= rva_out_reg_data_103_96_sva_dfm_4_mx0w0_3_0;
      rva_out_reg_data_111_104_sva_dfm_6_6_0 <= rva_out_reg_data_111_104_sva_dfm_4_mx0w0_6_0;
      rva_out_reg_data_119_112_sva_dfm_6_6_0 <= rva_out_reg_data_119_112_sva_dfm_4_mx0w0_6_0;
      rva_out_reg_data_95_88_sva_dfm_6_3_0 <= rva_out_reg_data_95_88_sva_dfm_7_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_base_input_and_tmp ) begin
      pe_manager_base_input_sva <= MUX_v_15_2_2(pe_manager_base_input_sva_dfm_3_1,
          while_if_while_if_and_2_nl, and_dcpl_220);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( (~((~((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6:4]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:7]!=3'b000))) & nor_721_cse
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:12]!=3'b000))) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]))
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & rva_in_PopNB_mioi_return_rsc_z_mxwt
        & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
        & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])))) & while_stage_0_3))
        & rva_in_reg_rw_and_5_cse ) begin
      pe_manager_base_input_sva_dfm_3_1 <= MUX_v_15_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[62:48]),
          pe_manager_base_input_sva_mx2, or_465_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_105_nl) & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_23_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_276_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_272_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_294_itm_1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_24_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_108_nl) & while_stage_0_5 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= MUX_s_1_2_2((pe_manager_base_weight_sva[0]), PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_3 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_45_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_27_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_195_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= rva_out_reg_data_30_25_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_196_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= rva_out_reg_data_23_17_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_197_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= rva_out_reg_data_15_9_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_198_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= rva_out_reg_data_35_32_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_199_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= rva_out_reg_data_39_36_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_200_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= rva_out_reg_data_46_40_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_201_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_4 <= rva_out_reg_data_62_56_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_202_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_4 <= rva_out_reg_data_55_48_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]))) & while_stage_0_4 )
        begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_29_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(reg_rva_in_reg_rw_sva_2_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= MUX_s_1_2_2(pe_manager_base_weight_sva_mx3_0, PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_46_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ reg_rva_in_reg_rw_sva_2_cse) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= input_read_req_valid_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_31_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= 6'b000000;
      rva_out_reg_data_23_17_sva_dfm_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_128_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= MUX_v_6_2_2(6'b000000, (pe_manager_base_weight_sva_mx2[14:9]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
      rva_out_reg_data_23_17_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_base_weight_sva_mx2[7:1]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_203_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= rva_out_reg_data_15_9_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_204_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= rva_out_reg_data_35_32_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_205_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= rva_out_reg_data_39_36_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_206_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= rva_out_reg_data_46_40_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_207_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_3 <= rva_out_reg_data_62_56_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_208_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_3 <= rva_out_reg_data_55_48_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= 1'b0;
      input_read_req_valid_lpi_1_dfm_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_35_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
      input_read_req_valid_lpi_1_dfm_1_2 <= input_read_req_valid_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_35_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_136_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= rva_out_reg_data_15_9_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_209_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= rva_out_reg_data_35_32_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_210_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= rva_out_reg_data_39_36_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_211_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= rva_out_reg_data_46_40_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_212_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_2 <= rva_out_reg_data_62_56_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_213_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_2 <= pe_config_input_counter_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (and_dcpl_479 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        & while_stage_0_3 ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_2_1,
          PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_479 & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1==4'b0100)
        & and_dcpl_488 & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2))
        & and_dcpl_212 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_1 <= 7'b0000000;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3;
      rva_out_reg_data_15_9_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_num_input_sva[7:1]),
          and_319_cse);
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_44_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= pe_config_is_cluster_sva;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1 <= pe_config_is_bias_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (or_dcpl_151 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
        | (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)))
        & and_dcpl_220 ) begin
      input_read_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_39_36_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_1_1 <= 7'b0000000;
      rva_out_reg_data_62_56_sva_dfm_1_1 <= 7'b0000000;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_143_cse ) begin
      rva_out_reg_data_35_32_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_6_nl
          & (signext_4_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1)) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_39_36_sva_dfm_1_1 <= (pe_manager_base_bias_sva[7:4]) & ({{3{and_319_cse}},
          and_319_cse}) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_46_40_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl
          & (signext_7_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1)) & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_62_56_sva_dfm_1_1 <= (pe_manager_base_input_sva_mx2[14:8])
          & ({{6{and_319_cse}}, and_319_cse}) & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_7_4 <= 4'b0000;
      weight_port_read_out_data_0_3_sva_dfm_1_3_0 <= 4'b0000;
      weight_port_read_out_data_0_1_sva_dfm_1_6_0 <= 7'b0000000;
    end
    else if ( and_1562_cse ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_7_4 <= MUX_v_4_2_2(4'b0000, mux1h_nl,
          not_2446_nl);
      weight_port_read_out_data_0_3_sva_dfm_1_3_0 <= MUX_v_4_2_2(4'b0000, mux1h_8_nl,
          not_2368_nl);
      weight_port_read_out_data_0_1_sva_dfm_1_6_0 <= MUX_v_7_2_2(7'b0000000, mux1h_11_nl,
          not_2449_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_5_4 <= 2'b00;
      weight_port_read_out_data_0_1_sva_dfm_1_7 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_1_7 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_1_6 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_131_ssc ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_5_4 <= MUX_v_2_2_2(2'b00, mux1h_9_nl,
          not_2448_nl);
      weight_port_read_out_data_0_1_sva_dfm_1_7 <= mux1h_2_nl & (~ or_dcpl);
      weight_port_read_out_data_0_2_sva_dfm_1_7 <= mux1h_1_nl & (~ or_dcpl_296);
      weight_port_read_out_data_0_2_sva_dfm_1_6 <= mux1h_15_nl & (~ or_dcpl_296);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_3_0 <= 4'b0000;
    end
    else if ( and_1568_tmp ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_3_0 <= MUX_v_4_2_2(4'b0000, mux1h_10_nl,
          not_2370_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1_6_0
          <= 7'b0000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1_6_0
          <= 7'b0000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_7_4
          <= 4'b0000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_3_0
          <= 4'b0000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_56_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_61_nl & (~ or_dcpl_300);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_86_nl,
          not_2357_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_66_nl & (~ or_dcpl_300);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_87_nl,
          not_2359_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_7_4
          <= MUX_v_4_2_2(4'b0000, weight_mem_banks_load_store_for_else_mux1h_71_nl,
          not_2360_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_3_0
          <= MUX_v_4_2_2(4'b0000, weight_mem_banks_load_store_for_else_mux1h_88_nl,
          not_2361_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_7_6
          <= 2'b00;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_5_0
          <= 6'b000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_68_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_7_6
          <= MUX_v_2_2_2(2'b00, weight_mem_banks_load_store_for_else_mux1h_76_nl,
          not_2362_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_5_0
          <= MUX_v_6_2_2(6'b000000, weight_mem_banks_load_store_for_else_mux1h_89_nl,
          not_2363_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_80_nl & (~ or_dcpl_300);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_90_nl,
          not_2365_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_75_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_7
          <= mux_493_nl & (~ and_dcpl_737);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, mux_494_nl, not_2367_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_225_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1 <= weight_port_read_out_data_0_0_sva_dfm_2_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_1 <= 2'b00;
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_0_1 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_0_0 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_185_ssc ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7 <= weight_port_read_out_data_0_0_sva_dfm_1_7;
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_0 <= weight_port_read_out_data_0_1_sva_dfm_1_7;
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_1 <= weight_port_read_out_data_0_2_sva_dfm_1_5_4;
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_0_1 <= weight_port_read_out_data_0_2_sva_dfm_1_7;
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_0_0 <= weight_port_read_out_data_0_2_sva_dfm_1_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_226_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0 <= weight_port_read_out_data_0_0_sva_dfm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_227_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_1 <= weight_port_read_out_data_0_1_sva_dfm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_2 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_228_enex5 ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_rsp_2 <= weight_port_read_out_data_0_2_sva_dfm_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_rsp_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_229_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_rsp_0 <= weight_port_read_out_data_0_3_sva_dfm_1_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_rsp_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_230_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_rsp_1 <= weight_port_read_out_data_0_3_sva_dfm_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_7 <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_1_6_0 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_189_ssc ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_7 <= weight_port_read_out_data_0_0_sva_dfm_mx0w0_7;
      weight_port_read_out_data_0_0_sva_dfm_1_6_0 <= MUX_v_7_2_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:9]),
          weight_port_read_out_data_0_0_sva_dfm_mx0w0_6_0, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_5_0 <=
          6'b000000;
    end
    else if ( weight_port_read_out_data_and_231_enex5 ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_5_0 <=
          reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_rsp_1
          <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_232_enex5 ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_rsp_1
          <= weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_5_rsp_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_233_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_5_rsp_0 <= weight_port_read_out_data_0_3_sva_dfm_4_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_5_rsp_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_234_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_5_rsp_1 <= weight_port_read_out_data_0_3_sva_dfm_4_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1_7_4 <= 4'b0000;
      weight_port_read_out_data_0_3_sva_dfm_1_1_3_0 <= 4'b0000;
    end
    else if ( and_1578_cse ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1_7_4 <= MUX1HOT_v_4_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001[7:4]),
          weight_port_read_out_data_0_3_sva_mx0_7_4, (weight_port_read_out_data_0_7_sva_dfm_mx0w2[7:4]),
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_nl,
          {and_dcpl_578 , and_dcpl_580 , and_dcpl_581 , and_dcpl_583});
      weight_port_read_out_data_0_3_sva_dfm_1_1_3_0 <= MUX1HOT_v_4_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000001[3:0]),
          weight_port_read_out_data_0_3_sva_mx0_3_0, (weight_port_read_out_data_0_7_sva_dfm_mx0w2[3:0]),
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_130_nl,
          {and_dcpl_578 , and_dcpl_580 , and_dcpl_581 , and_dcpl_583});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_7 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_1_1_6 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_1_1_5_4 <= 2'b00;
      weight_port_read_out_data_0_1_sva_dfm_1_1_7 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_130_ssc ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_7 <= MUX1HOT_s_1_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002[7]),
          weight_port_read_out_data_0_2_sva_mx0_7, weight_port_read_out_data_0_5_sva_dfm_mx0w2_7,
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_nl,
          {and_dcpl_578 , and_dcpl_580 , and_dcpl_581 , and_dcpl_583});
      weight_port_read_out_data_0_2_sva_dfm_1_1_6 <= MUX1HOT_s_1_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002[6]),
          weight_port_read_out_data_0_2_sva_mx0_6, (weight_port_read_out_data_0_5_sva_dfm_mx0w2_6_0[6]),
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_128_nl,
          {and_dcpl_578 , and_dcpl_580 , and_dcpl_581 , and_dcpl_583});
      weight_port_read_out_data_0_2_sva_dfm_1_1_5_4 <= MUX1HOT_v_2_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002[5:4]),
          weight_port_read_out_data_0_2_sva_mx0_5_4, (weight_port_read_out_data_0_5_sva_dfm_mx0w2_6_0[5:4]),
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_135_nl,
          {and_dcpl_578 , and_dcpl_580 , and_dcpl_581 , and_dcpl_583});
      weight_port_read_out_data_0_1_sva_dfm_1_1_7 <= MUX1HOT_s_1_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000[7]),
          weight_port_read_out_data_0_1_sva_mx0_7, weight_port_read_out_data_0_4_sva_dfm_mx0w2_7,
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_nl,
          {and_dcpl_578 , and_dcpl_580 , and_dcpl_581 , and_dcpl_583});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_3_0 <= 4'b0000;
    end
    else if ( mux_607_nl & PECoreRun_wen ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_3_0 <= MUX1HOT_v_4_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000002[3:0]),
          weight_port_read_out_data_0_2_sva_mx0_3_0, (weight_port_read_out_data_0_5_sva_dfm_mx0w2_6_0[3:0]),
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_136_nl,
          {and_dcpl_578 , and_dcpl_580 , and_dcpl_581 , and_dcpl_583});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_1_6_0 <= 7'b0000000;
    end
    else if ( mux_614_nl & PECoreRun_wen ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_1_6_0 <= MUX1HOT_v_7_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000000[6:0]),
          weight_port_read_out_data_0_1_sva_mx0_6_0, weight_port_read_out_data_0_4_sva_dfm_mx0w2_6_0,
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_129_nl,
          {and_dcpl_578 , and_dcpl_580 , and_dcpl_581 , and_dcpl_583});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (and_dcpl_41 | and_dcpl_33) ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7_1 <= MUX_s_1_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w0_7,
          weight_port_read_out_data_0_0_sva_dfm_3_7, and_dcpl_33);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0_1 <= 7'b0000000;
    end
    else if ( mux_617_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0_1 <= MUX_v_7_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w0_6_0,
          weight_port_read_out_data_0_0_sva_dfm_3_6_0, and_dcpl_33);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_5_0 <=
          6'b000000;
    end
    else if ( weight_port_read_out_data_and_235_enex5 ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_5_0 <=
          reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1[6:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_4_7_4 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_236_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_4_7_4 <= reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_4_3_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_237_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_4_3_0 <= reg_weight_port_read_out_data_0_3_sva_dfm_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_1_3 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_1_2_0 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_93_cse ) begin
      rva_out_reg_data_39_36_sva_dfm_4_1_3 <= MUX1HOT_s_1_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_3_0[3]),
          rva_out_reg_data_39_36_sva_dfm_6_mx1_3, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[39]),
          weight_port_read_out_data_0_4_sva_dfm_mx0w2_7, {PECore_PushAxiRsp_if_asn_89
          , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_39_36_sva_dfm_4_1_2_0 <= MUX1HOT_v_3_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_3_0[2:0]),
          rva_out_reg_data_39_36_sva_dfm_6_mx1_2_0, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[38:36]),
          (weight_port_read_out_data_0_4_sva_dfm_mx0w2_6_0[6:4]), {PECore_PushAxiRsp_if_asn_89
          , PECore_PushAxiRsp_if_asn_91 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_6_rsp_0 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_1 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_106_cse ) begin
      rva_out_reg_data_39_36_sva_dfm_6_rsp_0 <= rva_out_reg_data_39_36_sva_dfm_6_mx1_3;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_1 <= rva_out_reg_data_39_36_sva_dfm_6_mx1_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7
          <= 1'b0;
    end
    else if ( weight_mem_banks_load_store_for_else_and_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7
          <= MUX1HOT_s_1_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_nl,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000003[7]),
          weight_port_read_out_data_0_5_sva_mx0_7, {and_dcpl_583 , and_dcpl_655 ,
          and_dcpl_656});
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7
          <= MUX1HOT_s_1_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_nl,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7_0_s000004[7]),
          weight_port_read_out_data_0_4_sva_mx0_7, {and_dcpl_583 , and_dcpl_655 ,
          and_dcpl_656});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_87_80_sva_dfm_4_2_rsp_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_214_enex5 ) begin
      rva_out_reg_data_87_80_sva_dfm_4_2_rsp_1 <= rva_out_reg_data_87_80_sva_dfm_4_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_87_80_sva_dfm_6_7 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_6_7 <= 1'b0;
      rva_out_reg_data_111_104_sva_dfm_6_7 <= 1'b0;
      rva_out_reg_data_119_112_sva_dfm_6_7 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_6_6 <= 1'b0;
      rva_out_reg_data_95_88_sva_dfm_6_5_4 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_112_cse ) begin
      rva_out_reg_data_87_80_sva_dfm_6_7 <= MUX_s_1_2_2(rva_out_reg_data_87_80_sva_dfm_7_7,
          rva_out_reg_data_87_80_sva_dfm_8_7, while_asn_1039);
      rva_out_reg_data_95_88_sva_dfm_6_7 <= MUX_s_1_2_2(rva_out_reg_data_95_88_sva_dfm_7_7,
          rva_out_reg_data_95_88_sva_dfm_8_7, while_asn_1039);
      rva_out_reg_data_111_104_sva_dfm_6_7 <= MUX_s_1_2_2(rva_out_reg_data_111_104_sva_dfm_4_mx0w0_7,
          rva_out_reg_data_111_104_sva_dfm_7_7, while_asn_1039);
      rva_out_reg_data_119_112_sva_dfm_6_7 <= MUX_s_1_2_2(rva_out_reg_data_119_112_sva_dfm_4_mx0w0_7,
          rva_out_reg_data_119_112_sva_dfm_7_7, while_asn_1039);
      rva_out_reg_data_95_88_sva_dfm_6_6 <= MUX_s_1_2_2(rva_out_reg_data_95_88_sva_dfm_7_6,
          rva_out_reg_data_95_88_sva_dfm_8_6, while_asn_1039);
      rva_out_reg_data_95_88_sva_dfm_6_5_4 <= MUX_v_2_2_2(rva_out_reg_data_95_88_sva_dfm_7_5_4,
          rva_out_reg_data_95_88_sva_dfm_8_5_4, while_asn_1039);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_87_80_sva_dfm_4_5_rsp_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_215_enex5 ) begin
      rva_out_reg_data_87_80_sva_dfm_4_5_rsp_1 <= rva_out_reg_data_87_80_sva_dfm_4_4_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_87_80_sva_dfm_4_4_6_0 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_216_enex5 ) begin
      rva_out_reg_data_87_80_sva_dfm_4_4_6_0 <= reg_rva_out_reg_data_87_80_sva_dfm_4_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_3_rsp_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_217_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_103_96_sva_dfm_4_2_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_3_rsp_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_218_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_103_96_sva_dfm_4_2_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_219_enex5 ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_2 <= rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_119_112_sva_dfm_4_2_rsp_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_220_enex5 ) begin
      rva_out_reg_data_119_112_sva_dfm_4_2_rsp_1 <= rva_out_reg_data_119_112_sva_dfm_4_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_104_sva_dfm_4_2_rsp_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_221_enex5 ) begin
      rva_out_reg_data_111_104_sva_dfm_4_2_rsp_1 <= rva_out_reg_data_111_104_sva_dfm_4_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_2_7_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_222_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_2_7_4 <= rva_out_reg_data_103_96_sva_dfm_4_1_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_2_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_223_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_2_3_0 <= rva_out_reg_data_103_96_sva_dfm_4_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_224_enex5 ) begin
      rva_out_reg_data_95_88_sva_dfm_4_2_rsp_1_3_0 <= reg_rva_out_reg_data_95_88_sva_dfm_4_1_1_ftd_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_119_112_sva_dfm_4_5_rsp_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_225_enex5 ) begin
      rva_out_reg_data_119_112_sva_dfm_4_5_rsp_1 <= rva_out_reg_data_119_112_sva_dfm_4_4_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_104_sva_dfm_4_5_rsp_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_226_enex5 ) begin
      rva_out_reg_data_111_104_sva_dfm_4_5_rsp_1 <= rva_out_reg_data_111_104_sva_dfm_4_4_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_5_7_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_227_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_5_7_4 <= reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_4_5_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_228_enex5 ) begin
      rva_out_reg_data_103_96_sva_dfm_4_5_3_0 <= reg_rva_out_reg_data_103_96_sva_dfm_4_4_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_119_112_sva_dfm_4_4_6_0 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_229_enex5 ) begin
      rva_out_reg_data_119_112_sva_dfm_4_4_6_0 <= reg_rva_out_reg_data_119_112_sva_dfm_4_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_104_sva_dfm_4_4_6_0 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_230_enex5 ) begin
      rva_out_reg_data_111_104_sva_dfm_4_4_6_0 <= reg_rva_out_reg_data_111_104_sva_dfm_4_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_231_enex5 ) begin
      rva_out_reg_data_95_88_sva_dfm_4_5_rsp_1_rsp_2 <= rva_out_reg_data_95_88_sva_dfm_4_4_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_88_sva_dfm_4_4_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_232_enex5 ) begin
      rva_out_reg_data_95_88_sva_dfm_4_4_3_0 <= reg_rva_out_reg_data_95_88_sva_dfm_4_3_ftd_1_rsp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_159_enex5 | rva_out_reg_data_and_147_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_enexo <= rva_out_reg_data_and_159_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_158_enex5 | rva_out_reg_data_and_148_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_enexo <= rva_out_reg_data_and_158_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_157_enex5 | rva_out_reg_data_and_149_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_7_enexo <= rva_out_reg_data_and_157_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_164_enex5 | rva_out_reg_data_and_150_enex5 ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_4_enexo <= rva_out_reg_data_and_164_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_167_enex5 | rva_out_reg_data_and_151_enex5 ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_4_enexo <= rva_out_reg_data_and_167_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_168_enex5 | rva_out_reg_data_and_152_enex5 ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_4_enexo <= rva_out_reg_data_and_168_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_162_enex5 | rva_out_reg_data_and_153_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_4_enexo <= rva_out_reg_data_and_162_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_160_enex5 | rva_out_reg_data_and_154_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo <= rva_out_reg_data_and_160_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_163_enex5 | rva_out_reg_data_and_155_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_enexo <= rva_out_reg_data_and_163_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_161_enex5 | rva_out_reg_data_and_156_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo <= rva_out_reg_data_and_161_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_51_enex5 | input_mem_banks_read_read_data_and_47_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo
          <= input_mem_banks_read_read_data_and_51_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_52_enex5 | input_mem_banks_read_read_data_and_48_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo
          <= input_mem_banks_read_read_data_and_52_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_53_enex5 | input_mem_banks_read_read_data_and_49_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo
          <= input_mem_banks_read_read_data_and_53_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_54_enex5 | input_mem_banks_read_read_data_and_50_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo
          <= input_mem_banks_read_read_data_and_54_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_16_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1446_cse | act_port_reg_data_and_19_enex5 ) begin
      reg_act_port_reg_data_16_0_sva_dfm_1_1_enexo <= and_1446_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_240_224_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1446_cse | act_port_reg_data_and_20_enex5 ) begin
      reg_act_port_reg_data_240_224_sva_dfm_1_1_enexo <= and_1446_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_208_192_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1446_cse | act_port_reg_data_and_21_enex5 ) begin
      reg_act_port_reg_data_208_192_sva_dfm_1_1_enexo <= and_1446_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_176_160_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1446_cse | act_port_reg_data_and_22_enex5 ) begin
      reg_act_port_reg_data_176_160_sva_dfm_1_1_enexo <= and_1446_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_1_enex5 | input_mem_banks_read_1_read_data_and_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_1_read_data_and_1_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp | weight_port_read_out_data_and_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= data_in_tmp_operator_2_for_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_190_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_191_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_192_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_193_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_194_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_195_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_196_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_197_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_198_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_199_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_200_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_201_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_202_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_203_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_204_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_205_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_206_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000001
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_207_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000002
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_208_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000003
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_209_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000004
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_210_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000005
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_211_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000006
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_212_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000007
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_213_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000008
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_214_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000009
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_215_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000010
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_216_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000011
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_217_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000012
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_218_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000013
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_219_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000014
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_31_tmp | weight_port_read_out_data_and_31_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_8_7000000
          <= data_in_tmp_operator_2_for_and_31_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_2_enex5 | input_mem_banks_read_1_read_data_and_1_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= input_mem_banks_read_1_read_data_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( weight_read_addrs_and_7_cse | weight_read_addrs_and_28_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= weight_read_addrs_and_7_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_enexo <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo
          <= 1'b1;
    end
    else if ( PECoreRun_wen | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo
          <= PECoreRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= 1'b1;
    end
    else if ( weight_read_addrs_and_7_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= weight_read_addrs_and_7_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_enexo_1 <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_enexo_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo_1
          <= 1'b1;
    end
    else if ( PECoreRun_wen | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 )
        begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo_1
          <= PECoreRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= 1'b1;
    end
    else if ( weight_read_addrs_and_7_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= weight_read_addrs_and_7_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= 1'b1;
    end
    else if ( operator_15_false_1_and_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= operator_15_false_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_64_enex5 | weight_write_data_data_and_48_enex5
        ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_64_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_65_enex5 | weight_write_data_data_and_49_enex5
        ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_65_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_66_enex5 | weight_write_data_data_and_50_enex5
        ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_67_enex5 | weight_write_data_data_and_51_enex5
        ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_68_enex5 | weight_write_data_data_and_52_enex5
        ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_69_enex5 | weight_write_data_data_and_53_enex5
        ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_70_enex5 | weight_write_data_data_and_54_enex5
        ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_70_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_71_enex5 | weight_write_data_data_and_55_enex5
        ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_71_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_72_enex5 | weight_write_data_data_and_56_enex5
        ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_72_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_73_enex5 | weight_write_data_data_and_57_enex5
        ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_73_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_74_enex5 | weight_write_data_data_and_58_enex5
        ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_74_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_75_enex5 | weight_write_data_data_and_59_enex5
        ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_75_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_76_enex5 | weight_write_data_data_and_60_enex5
        ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_76_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_77_enex5 | weight_write_data_data_and_61_enex5
        ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_77_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_78_enex5 | weight_write_data_data_and_62_enex5
        ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_78_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_79_enex5 | weight_write_data_data_and_63_enex5
        ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_79_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_write_addrs_and_2_enex5 | weight_write_addrs_and_enex5 ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= weight_write_addrs_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_64_enex5 ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_65_enex5 ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_66_enex5 ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_67_enex5 ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_68_enex5 ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_69_enex5 ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_70_enex5 ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_71_enex5 ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_72_enex5 ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_73_enex5 ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_74_enex5 ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_75_enex5 ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_76_enex5 ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_77_enex5 ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_78_enex5 ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_79_enex5 ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_input_enexo <= 1'b1;
    end
    else if ( pe_manager_base_input_and_tmp | weight_write_addrs_and_2_enex5 ) begin
      reg_pe_manager_base_input_enexo <= pe_manager_base_input_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_read_addrs_and_29_enex5 ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_config_num_output_enexo <= 1'b1;
    end
    else if ( pe_config_num_manager_and_cse | pe_config_UpdateManagerCounter_if_if_and_enex5
        ) begin
      reg_pe_config_num_output_enexo <= pe_config_num_manager_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_read_addrs_and_30_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_data_sva_1_enexo <= 1'b1;
    end
    else if ( rva_in_reg_data_and_tmp | PEManager_15U_PEManagerWrite_and_enex5 )
        begin
      reg_rva_in_reg_data_sva_1_enexo <= rva_in_reg_data_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_225_enex5 | weight_port_read_out_data_and_220_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_225_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_55_enex5 | input_mem_banks_read_read_data_and_51_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo
          <= input_mem_banks_read_read_data_and_55_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_56_enex5 | input_mem_banks_read_read_data_and_52_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo
          <= input_mem_banks_read_read_data_and_56_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_57_enex5 | input_mem_banks_read_read_data_and_53_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo
          <= input_mem_banks_read_read_data_and_57_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_58_enex5 | input_mem_banks_read_read_data_and_54_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo
          <= input_mem_banks_read_read_data_and_58_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 | input_mem_banks_read_1_read_data_and_2_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_1_read_data_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_169_enex5 | rva_out_reg_data_and_157_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= rva_out_reg_data_and_169_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_170_enex5 | rva_out_reg_data_and_158_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= rva_out_reg_data_and_170_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_171_enex5 | rva_out_reg_data_and_159_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= rva_out_reg_data_and_171_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_172_enex5 | rva_out_reg_data_and_160_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= rva_out_reg_data_and_172_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_173_enex5 | rva_out_reg_data_and_161_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo <= rva_out_reg_data_and_173_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_174_enex5 | rva_out_reg_data_and_162_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo <= rva_out_reg_data_and_174_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_175_enex5 | rva_out_reg_data_and_163_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo <= rva_out_reg_data_and_175_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_176_enex5 | rva_out_reg_data_and_164_enex5 ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_3_enexo <= rva_out_reg_data_and_176_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_217_enex5 | rva_out_reg_data_and_165_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_3_enexo <= rva_out_reg_data_and_217_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_218_enex5 | rva_out_reg_data_and_166_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_218_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_180_enex5 | rva_out_reg_data_and_167_enex5 ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_3_enexo <= rva_out_reg_data_and_180_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_181_enex5 | rva_out_reg_data_and_168_enex5 ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_3_enexo <= rva_out_reg_data_and_181_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_227_enex5 | weight_port_read_out_data_and_221_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_227_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_228_enex5 | weight_port_read_out_data_and_222_enex5
        ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo <= weight_port_read_out_data_and_228_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= 1'b1;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_1_for_and_cse | weight_mem_write_arbxbar_xbar_for_empty_and_enex5
        ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= weight_mem_write_arbxbar_xbar_for_1_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_59_enex5 | input_mem_banks_read_read_data_and_55_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= input_mem_banks_read_read_data_and_59_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_60_enex5 | input_mem_banks_read_read_data_and_56_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= input_mem_banks_read_read_data_and_60_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_61_enex5 | input_mem_banks_read_read_data_and_57_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= input_mem_banks_read_read_data_and_61_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_62_enex5 | input_mem_banks_read_read_data_and_58_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= input_mem_banks_read_read_data_and_62_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp | input_mem_banks_read_1_read_data_and_3_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= input_mem_banks_read_1_read_data_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_182_enex5 | rva_out_reg_data_and_169_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= rva_out_reg_data_and_182_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_183_enex5 | rva_out_reg_data_and_170_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= rva_out_reg_data_and_183_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_184_enex5 | rva_out_reg_data_and_171_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= rva_out_reg_data_and_184_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_229_enex5 | weight_port_read_out_data_and_223_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_enexo <= weight_port_read_out_data_and_229_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_230_enex5 | weight_port_read_out_data_and_224_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_230_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_185_enex5 | rva_out_reg_data_and_172_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= rva_out_reg_data_and_185_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_186_enex5 | rva_out_reg_data_and_173_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo <= rva_out_reg_data_and_186_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_187_enex5 | rva_out_reg_data_and_174_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo <= rva_out_reg_data_and_187_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_188_enex5 | rva_out_reg_data_and_175_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo <= rva_out_reg_data_and_188_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_189_enex5 | rva_out_reg_data_and_176_enex5 ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_2_enexo <= rva_out_reg_data_and_189_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_220_enex5 | rva_out_reg_data_and_177_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_220_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_221_enex5 | rva_out_reg_data_and_178_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_221_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_214_enex5 | rva_out_reg_data_and_179_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_214_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_190_enex5 | rva_out_reg_data_and_180_enex5 ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_2_enexo <= rva_out_reg_data_and_190_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_191_enex5 | rva_out_reg_data_and_181_enex5 ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_2_enexo <= rva_out_reg_data_and_191_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_63_enex5 | input_mem_banks_read_read_data_and_59_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= input_mem_banks_read_read_data_and_63_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_189_ssc | input_mem_banks_read_read_data_and_60_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo <= weight_port_read_out_data_and_189_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_64_enex5 | input_mem_banks_read_read_data_and_61_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= input_mem_banks_read_read_data_and_64_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_65_enex5 | input_mem_banks_read_read_data_and_62_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= input_mem_banks_read_read_data_and_65_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_192_enex5 | rva_out_reg_data_and_182_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_4_enexo <= rva_out_reg_data_and_192_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_193_enex5 | rva_out_reg_data_and_183_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_4_enexo <= rva_out_reg_data_and_193_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_194_enex5 | rva_out_reg_data_and_184_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_6_enexo <= rva_out_reg_data_and_194_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1489_cse | rva_out_reg_data_and_185_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= and_1489_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1489_cse | rva_out_reg_data_and_186_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo <= and_1489_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1489_cse | rva_out_reg_data_and_187_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo <= and_1489_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1489_cse | rva_out_reg_data_and_188_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo <= and_1489_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_98_cse | rva_out_reg_data_and_189_enex5 ) begin
      reg_rva_out_reg_data_127_120_sva_dfm_4_1_enexo <= rva_out_reg_data_and_98_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( input_read_req_valid_and_4_cse | rva_out_reg_data_and_190_enex5 ) begin
      reg_rva_out_reg_data_79_72_sva_dfm_4_1_enexo <= input_read_req_valid_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( input_read_req_valid_and_4_cse | rva_out_reg_data_and_191_enex5 ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_4_1_enexo <= input_read_req_valid_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_44_tmp | input_mem_banks_read_read_data_and_63_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_read_data_and_44_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_44_tmp | input_mem_banks_read_read_data_and_64_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1 <= input_mem_banks_read_read_data_and_44_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_44_tmp | input_mem_banks_read_read_data_and_65_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2 <= input_mem_banks_read_read_data_and_44_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( weight_mem_banks_load_store_for_else_and_68_ssc | rva_out_reg_data_and_192_enex5
        ) begin
      reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_1_enexo
          <= weight_mem_banks_load_store_for_else_and_68_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( weight_mem_banks_load_store_for_else_and_68_ssc | rva_out_reg_data_and_193_enex5
        ) begin
      reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_1_enexo
          <= weight_mem_banks_load_store_for_else_and_68_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( weight_mem_banks_load_store_for_else_and_75_ssc | rva_out_reg_data_and_194_enex5
        ) begin
      reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1_1_enexo
          <= weight_mem_banks_load_store_for_else_and_75_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_46_enex5 | input_mem_banks_read_read_data_and_45_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_read_data_and_46_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_128_cse | rva_out_reg_data_and_195_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= rva_out_reg_data_and_128_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_128_cse | rva_out_reg_data_and_196_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= rva_out_reg_data_and_128_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_203_enex5 | rva_out_reg_data_and_197_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= rva_out_reg_data_and_203_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_204_enex5 | rva_out_reg_data_and_198_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= rva_out_reg_data_and_204_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_205_enex5 | rva_out_reg_data_and_199_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= rva_out_reg_data_and_205_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_206_enex5 | rva_out_reg_data_and_200_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= rva_out_reg_data_and_206_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_207_enex5 | rva_out_reg_data_and_201_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo <= rva_out_reg_data_and_207_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_208_enex5 | rva_out_reg_data_and_202_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo <= rva_out_reg_data_and_208_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp | input_mem_banks_read_read_data_and_46_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1 <= input_mem_banks_read_1_read_data_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_136_enex5 | rva_out_reg_data_and_203_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= rva_out_reg_data_and_136_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_209_enex5 | rva_out_reg_data_and_204_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= rva_out_reg_data_and_209_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_210_enex5 | rva_out_reg_data_and_205_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= rva_out_reg_data_and_210_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_211_enex5 | rva_out_reg_data_and_206_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= rva_out_reg_data_and_211_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_212_enex5 | rva_out_reg_data_and_207_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo <= rva_out_reg_data_and_212_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_213_enex5 | rva_out_reg_data_and_208_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo <= rva_out_reg_data_and_213_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse | rva_out_reg_data_and_136_enex5
        ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_42_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_143_cse | rva_out_reg_data_and_209_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= rva_out_reg_data_and_143_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_143_cse | rva_out_reg_data_and_210_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= rva_out_reg_data_and_143_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_143_cse | rva_out_reg_data_and_211_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= rva_out_reg_data_and_143_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_143_cse | rva_out_reg_data_and_212_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo <= rva_out_reg_data_and_143_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_config_input_counter_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( and_1441_tmp | rva_out_reg_data_and_213_enex5 ) begin
      reg_pe_config_input_counter_sva_dfm_1_enexo <= and_1441_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_226_enex5 | weight_port_read_out_data_and_225_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_226_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo_1 <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_189_ssc | weight_port_read_out_data_and_226_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo_1 <= weight_port_read_out_data_and_189_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1562_cse | weight_port_read_out_data_and_227_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo <= and_1562_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( and_1568_tmp | weight_port_read_out_data_and_228_enex5 ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_1_2_enexo <= and_1568_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( and_1562_cse | weight_port_read_out_data_and_229_enex5 ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_enexo <= and_1562_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1562_cse | weight_port_read_out_data_and_230_enex5 ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_1_enexo <= and_1562_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_220_enex5 | weight_port_read_out_data_and_231_enex5
        ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_1_enexo
          <= weight_port_read_out_data_and_220_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_235_enex5 | weight_port_read_out_data_and_232_enex5
        ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_1_enexo
          <= weight_port_read_out_data_and_235_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_236_enex5 | weight_port_read_out_data_and_233_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_enexo <= weight_port_read_out_data_and_236_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_237_enex5 | weight_port_read_out_data_and_234_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_1_enexo <= weight_port_read_out_data_and_237_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_221_enex5 | weight_port_read_out_data_and_235_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_221_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_223_enex5 | weight_port_read_out_data_and_236_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_enexo <= weight_port_read_out_data_and_223_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_224_enex5 | weight_port_read_out_data_and_237_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_224_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( input_read_req_valid_and_4_cse | rva_out_reg_data_and_214_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_1_1_enexo <= input_read_req_valid_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_216_enex5 | rva_out_reg_data_and_215_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_4_1_enexo <= rva_out_reg_data_and_216_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_179_enex5 | rva_out_reg_data_and_216_enex5 ) begin
      reg_rva_out_reg_data_87_80_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_179_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_222_enex5 | rva_out_reg_data_and_217_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_2_enexo <= rva_out_reg_data_and_222_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_223_enex5 | rva_out_reg_data_and_218_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_223_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_2_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_224_enex5 | rva_out_reg_data_and_219_enex5 ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_2_3_enexo <= rva_out_reg_data_and_224_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_98_cse | rva_out_reg_data_and_220_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_1_1_enexo <= rva_out_reg_data_and_98_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_98_cse | rva_out_reg_data_and_221_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_1_1_enexo <= rva_out_reg_data_and_98_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_98_cse | rva_out_reg_data_and_222_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_1_enexo <= rva_out_reg_data_and_98_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_98_cse | rva_out_reg_data_and_223_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_1_1_enexo <= rva_out_reg_data_and_98_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_3_enexo <= 1'b1;
    end
    else if ( input_read_req_valid_and_4_cse | rva_out_reg_data_and_224_enex5 ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_1_3_enexo <= input_read_req_valid_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_229_enex5 | rva_out_reg_data_and_225_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_4_1_enexo <= rva_out_reg_data_and_229_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_230_enex5 | rva_out_reg_data_and_226_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_4_1_enexo <= rva_out_reg_data_and_230_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_165_enex5 | rva_out_reg_data_and_227_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_enexo <= rva_out_reg_data_and_165_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_166_enex5 | rva_out_reg_data_and_228_enex5 ) begin
      reg_rva_out_reg_data_103_96_sva_dfm_4_4_1_enexo <= rva_out_reg_data_and_166_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_177_enex5 | rva_out_reg_data_and_229_enex5 ) begin
      reg_rva_out_reg_data_119_112_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_177_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_178_enex5 | rva_out_reg_data_and_230_enex5 ) begin
      reg_rva_out_reg_data_111_104_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_178_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_232_enex5 | rva_out_reg_data_and_231_enex5 ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_4_3_enexo <= rva_out_reg_data_and_232_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_219_enex5 | rva_out_reg_data_and_232_enex5 ) begin
      reg_rva_out_reg_data_95_88_sva_dfm_4_3_3_enexo <= rva_out_reg_data_and_219_enex5;
    end
  end
  assign nl_operator_4_false_acc_nl = pe_config_manager_counter_sva_mx1 + 4'b0001;
  assign operator_4_false_acc_nl = nl_operator_4_false_acc_nl[3:0];
  assign pe_config_UpdateManagerCounter_if_not_7_nl = ~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  assign nl_input_read_addrs_sva_1_1  = pe_config_input_counter_sva_mx1 + pe_manager_base_input_sva_mx1_7_0;
  assign PECore_RunScale_if_for_2_scaled_val_mul_1_nl = (accum_vector_data_1_19_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_3_scaled_val_mul_1_nl = (accum_vector_data_2_19_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_4_scaled_val_mul_1_nl = (accum_vector_data_3_19_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_5_scaled_val_mul_1_nl = (accum_vector_data_4_19_0_sva)
      * 8'b10100111;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_119_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_1_nl = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:120]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:120]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:120]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:120]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_8_mx0[119:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_238_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_248_itm_1});
  assign mux_7_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_7_lpi_1_dfm_1, (~ rva_in_reg_rw_sva_4),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_10_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_6_lpi_1_dfm_1, (~ rva_in_reg_rw_sva_st_1_4),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_136_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_134_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_151_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_188_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_28_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign nor_692_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ or_tmp_586));
  assign mux_538_nl = MUX_s_1_2_2(or_tmp_586, nor_692_nl, while_stage_0_6);
  assign mux_539_nl = MUX_s_1_2_2(mux_538_nl, or_tmp_586, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_48_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[7:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl);
  assign nor_483_nl = ~((~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_11_nl = MUX_s_1_2_2(nor_483_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_138_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_80_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[7:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_138_nl);
  assign nor_484_nl = ~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_12_nl = MUX_s_1_2_2(nor_484_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_38_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign or_37_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | and_797_cse
      | and_798_cse | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign mux_14_nl = MUX_s_1_2_2(or_37_nl, or_tmp_19, weight_mem_read_arbxbar_arbiters_next_7_3_sva);
  assign mux_15_nl = MUX_s_1_2_2(or_38_nl, mux_14_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign or_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])) | weight_mem_read_arbxbar_arbiters_next_7_6_sva
      | (~ weight_mem_read_arbxbar_arbiters_next_7_3_sva) | or_tmp_19;
  assign mux_16_nl = MUX_s_1_2_2(mux_15_nl, or_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign or_39_nl = (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ mux_16_nl);
  assign or_31_nl = (~(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3))
      | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_13_nl = MUX_s_1_2_2(or_31_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3,
      or_tmp_14);
  assign mux_17_nl = MUX_s_1_2_2(or_39_nl, mux_13_nl, while_stage_0_5);
  assign or_28_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_18_nl = MUX_s_1_2_2(mux_17_nl, or_28_nl, while_stage_0_6);
  assign or_53_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign or_52_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])
      | and_799_cse | and_800_cse | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign mux_20_nl = MUX_s_1_2_2(or_52_nl, or_tmp_32, weight_mem_read_arbxbar_arbiters_next_6_3_sva);
  assign mux_21_nl = MUX_s_1_2_2(or_53_nl, mux_20_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign or_48_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])) | (~
      weight_mem_read_arbxbar_arbiters_next_6_3_sva) | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | or_tmp_32;
  assign mux_22_nl = MUX_s_1_2_2(mux_21_nl, or_48_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_54_nl = (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ mux_22_nl);
  assign or_43_nl = (~(Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6 |
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3)) | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_19_nl = MUX_s_1_2_2(or_43_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3,
      or_tmp_26);
  assign mux_23_nl = MUX_s_1_2_2(or_54_nl, mux_19_nl, while_stage_0_5);
  assign or_40_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_24_nl = MUX_s_1_2_2(mux_23_nl, or_40_nl, while_stage_0_6);
  assign mux_25_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_3, (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign nor_693_nl = ~((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign nor_694_nl = ~((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | (~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | (~ reg_rva_in_reg_rw_sva_st_1_1_cse));
  assign mux_540_nl = MUX_s_1_2_2(nor_693_nl, nor_694_nl, while_stage_0_3);
  assign mux_541_nl = MUX_s_1_2_2(mux_540_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2,
      while_stage_0_4);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl
      = MUX_v_11_2_2(11'b00000000000, PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl
      = MUX_v_4_2_2(4'b0000, pe_config_manager_counter_sva_mx1, PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign and_662_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & reg_rva_in_PopNB_mioi_iswt0_cse & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))
      & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl = (state_mux_1_cse!=2'b00)
      | state_0_sva_mx1;
  assign PECore_UpdateFSM_switch_lp_or_nl = PECore_UpdateFSM_switch_lp_equal_tmp_6
      | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  assign PECore_UpdateFSM_switch_lp_mux1h_15_nl = MUX1HOT_v_2_3_2((signext_2_1(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl)),
      2'b01, 2'b10, {PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      , PECore_UpdateFSM_switch_lp_or_nl , PECore_RunScale_PECore_RunScale_if_and_1_svs_1});
  assign PECore_UpdateFSM_switch_lp_nor_8_nl = ~(PECore_PushOutput_PECore_PushOutput_if_and_svs_1
      | PECore_UpdateFSM_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_and_1_nl = MUX_v_2_2_2(2'b00, PECore_UpdateFSM_switch_lp_mux1h_15_nl,
      PECore_UpdateFSM_switch_lp_nor_8_nl);
  assign nor_705_nl = ~((~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1);
  assign mux_542_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_3_1, nor_705_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nand_73_nl = ~(PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign or_1015_nl = (~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
  assign mux_543_nl = MUX_s_1_2_2(nand_73_nl, or_1015_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nl_operator_8_false_acc_sdt_sva_1  = conv_u2s_8_9(pe_config_num_output_sva)
      + 9'b111111111;
  assign nl_ProductSum_for_acc_39_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_32_z)
      + conv_u2u_18_20({Datapath_for_2_ProductSum_for_acc_2_1_17 , Datapath_for_2_ProductSum_for_acc_2_1_16_0})
      + conv_u2u_18_20({Datapath_for_2_ProductSum_for_acc_3_1_17 , Datapath_for_2_ProductSum_for_acc_3_1_16_0});
  assign ProductSum_for_acc_39_nl = nl_ProductSum_for_acc_39_nl[19:0];
  assign nl_ProductSum_for_acc_38_nl = ProductSum_for_acc_39_nl + ProductSum_for_acc_40_itm_1
      + conv_u2s_19_20(ProductSum_for_acc_41_itm_1);
  assign ProductSum_for_acc_38_nl = nl_ProductSum_for_acc_38_nl[19:0];
  assign PECore_UpdateFSM_switch_lp_not_21_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_31_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_48_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_47_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_46_z);
  assign ProductSum_for_acc_31_nl = nl_ProductSum_for_acc_31_nl[19:0];
  assign nl_ProductSum_for_acc_32_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_45_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_44_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_43_z);
  assign ProductSum_for_acc_32_nl = nl_ProductSum_for_acc_32_nl[19:0];
  assign nl_ProductSum_for_acc_33_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_42_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_41_z);
  assign ProductSum_for_acc_33_nl = nl_ProductSum_for_acc_33_nl[18:0];
  assign nl_ProductSum_for_acc_30_nl = ProductSum_for_acc_31_nl + ProductSum_for_acc_32_nl
      + conv_u2s_19_20(ProductSum_for_acc_33_nl);
  assign ProductSum_for_acc_30_nl = nl_ProductSum_for_acc_30_nl[19:0];
  assign PECore_UpdateFSM_switch_lp_not_36_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_27_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_56_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_55_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_54_z);
  assign ProductSum_for_acc_27_nl = nl_ProductSum_for_acc_27_nl[19:0];
  assign nl_ProductSum_for_acc_28_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_53_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_52_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_51_z);
  assign ProductSum_for_acc_28_nl = nl_ProductSum_for_acc_28_nl[19:0];
  assign nl_ProductSum_for_acc_29_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_50_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_49_z);
  assign ProductSum_for_acc_29_nl = nl_ProductSum_for_acc_29_nl[18:0];
  assign nl_ProductSum_for_acc_26_nl = ProductSum_for_acc_27_nl + ProductSum_for_acc_28_nl
      + conv_u2s_19_20(ProductSum_for_acc_29_nl);
  assign ProductSum_for_acc_26_nl = nl_ProductSum_for_acc_26_nl[19:0];
  assign PECore_UpdateFSM_switch_lp_not_34_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_23_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_z)
      + conv_u2u_18_20({Datapath_for_4_ProductSum_for_acc_2_1_17 , Datapath_for_4_ProductSum_for_acc_2_1_16_0})
      + conv_u2u_18_20({Datapath_for_4_ProductSum_for_acc_3_1_17 , Datapath_for_4_ProductSum_for_acc_3_1_16_0});
  assign ProductSum_for_acc_23_nl = nl_ProductSum_for_acc_23_nl[19:0];
  assign nl_ProductSum_for_acc_22_nl = ProductSum_for_acc_23_nl + ProductSum_for_acc_24_itm_1
      + conv_u2s_19_20(ProductSum_for_acc_25_itm_1);
  assign ProductSum_for_acc_22_nl = nl_ProductSum_for_acc_22_nl[19:0];
  assign PECore_UpdateFSM_switch_lp_not_35_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_234_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[127:120]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_234_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_278_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_138_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[118:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_278_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_277_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_137_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[110:104]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_277_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_249_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_174_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_189_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_204_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_219_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_250_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_175_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_190_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_205_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_220_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_251_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_176_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_191_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_206_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_221_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_252_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_177_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_192_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_207_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_222_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_253_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_178_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_193_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_208_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_223_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_254_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_179_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_194_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_209_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_224_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_240_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_255_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_180_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_195_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_210_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_225_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_241_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_181_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_196_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_211_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_226_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_242_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_257_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_182_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_197_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_212_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_227_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_243_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_244_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_246_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign and_1171_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])
      & (~ or_dcpl_298);
  assign and_1172_nl = and_dcpl_657 & (~ or_dcpl_298);
  assign and_1173_nl = nor_436_cse & (~ or_dcpl_298);
  assign mux1h_3_nl = MUX1HOT_v_8_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[63:56]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[63:56]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[63:56]),
      {and_1171_nl , and_1172_nl , and_1173_nl});
  assign not_2374_nl = ~ or_dcpl_298;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_198_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_201_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_202_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_203_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_228_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_229_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_231_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_233_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_199_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_200_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_245_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_140_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_230_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_232_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign or_222_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1;
  assign mux_40_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_5_lpi_1_dfm_1, or_222_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_221_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_itm_1;
  assign mux_39_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_5_lpi_1_dfm_1, or_221_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_41_nl = MUX_s_1_2_2(mux_40_nl, mux_39_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign or_220_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_5_lpi_1_dfm_1;
  assign mux_42_nl = MUX_s_1_2_2(mux_41_nl, or_220_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp);
  assign or_236_nl = (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])))
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign or_234_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 | and_801_cse));
  assign mux_43_nl = MUX_s_1_2_2(or_236_nl, or_234_nl, while_stage_0_5);
  assign or_241_nl = (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4])))
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign or_239_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 | and_802_cse));
  assign mux_44_nl = MUX_s_1_2_2(or_241_nl, or_239_nl, while_stage_0_5);
  assign or_253_nl = (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_15_tmp))
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign or_251_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_15_tmp)) |
      (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign mux_54_nl = MUX_s_1_2_2(or_253_nl, or_251_nl, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign or_249_nl = (~(weight_mem_read_arbxbar_arbiters_next_3_5_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]))
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_15_tmp)) |
      (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign mux_55_nl = MUX_s_1_2_2(mux_54_nl, or_249_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign mux_53_nl = MUX_s_1_2_2(or_tmp_75, or_dcpl_75, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1);
  assign mux_56_nl = MUX_s_1_2_2(mux_55_nl, mux_53_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign mux_655_nl = MUX_s_1_2_2(or_tmp_75, or_dcpl_75, and_770_cse);
  assign mux_52_nl = MUX_s_1_2_2(mux_655_nl, or_dcpl_75, weight_mem_read_arbxbar_arbiters_next_3_2_sva);
  assign mux_57_nl = MUX_s_1_2_2(mux_56_nl, mux_52_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign mux_657_nl = MUX_s_1_2_2(or_tmp_75, or_dcpl_75, and_770_cse);
  assign mux_474_nl = MUX_s_1_2_2(mux_657_nl, or_dcpl_75, and_776_cse);
  assign mux_51_nl = MUX_s_1_2_2(mux_474_nl, or_dcpl_75, weight_mem_read_arbxbar_arbiters_next_3_6_sva);
  assign mux_58_nl = MUX_s_1_2_2(mux_57_nl, mux_51_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign mux_659_nl = MUX_s_1_2_2(or_tmp_75, or_dcpl_75, and_770_cse);
  assign mux_468_nl = MUX_s_1_2_2(mux_659_nl, or_dcpl_75, and_776_cse);
  assign mux_47_nl = MUX_s_1_2_2(mux_468_nl, or_dcpl_75, and_771_cse);
  assign mux_50_nl = MUX_s_1_2_2(mux_47_nl, or_dcpl_75, weight_mem_read_arbxbar_arbiters_next_3_3_sva);
  assign mux_59_nl = MUX_s_1_2_2(mux_58_nl, mux_50_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign mux_505_nl = MUX_s_1_2_2(or_tmp_75, or_dcpl_75, and_770_cse);
  assign mux_46_nl = MUX_s_1_2_2(mux_505_nl, or_dcpl_75, and_776_cse);
  assign mux_464_nl = MUX_s_1_2_2(mux_46_nl, or_dcpl_75, and_771_cse);
  assign mux_48_nl = MUX_s_1_2_2(mux_464_nl, or_dcpl_75, and_773_cse);
  assign mux_49_nl = MUX_s_1_2_2(mux_48_nl, or_dcpl_75, weight_mem_read_arbxbar_arbiters_next_3_1_sva);
  assign mux_60_nl = MUX_s_1_2_2(mux_59_nl, mux_49_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign or_244_nl = (~(and_774_cse | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1))
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_61_nl = MUX_s_1_2_2(mux_60_nl, or_244_nl, while_stage_0_5);
  assign or_262_nl = (~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp)
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign or_261_nl = (~(weight_mem_read_arbxbar_arbiters_next_2_5_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]))
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_11_tmp)) |
      (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign mux_73_nl = MUX_s_1_2_2(or_262_nl, or_261_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign mux_72_nl = MUX_s_1_2_2(or_tmp_87, or_dcpl_75, weight_mem_read_arbxbar_arbiters_next_2_4_sva);
  assign mux_74_nl = MUX_s_1_2_2(mux_73_nl, mux_72_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign mux_656_nl = MUX_s_1_2_2(or_tmp_87, or_dcpl_75, and_766_cse);
  assign mux_71_nl = MUX_s_1_2_2(mux_656_nl, or_dcpl_75, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1);
  assign mux_75_nl = MUX_s_1_2_2(mux_74_nl, mux_71_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign mux_658_nl = MUX_s_1_2_2(or_tmp_87, or_dcpl_75, and_766_cse);
  assign mux_63_nl = MUX_s_1_2_2(mux_658_nl, or_dcpl_75, and_740_cse);
  assign mux_70_nl = MUX_s_1_2_2(mux_63_nl, or_dcpl_75, weight_mem_read_arbxbar_arbiters_next_2_3_sva);
  assign mux_76_nl = MUX_s_1_2_2(mux_75_nl, mux_70_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign mux_660_nl = MUX_s_1_2_2(or_tmp_87, or_dcpl_75, and_766_cse);
  assign mux_470_nl = MUX_s_1_2_2(mux_660_nl, or_dcpl_75, and_740_cse);
  assign mux_64_nl = MUX_s_1_2_2(mux_470_nl, or_dcpl_75, and_767_cse);
  assign mux_69_nl = MUX_s_1_2_2(mux_64_nl, or_dcpl_75, weight_mem_read_arbxbar_arbiters_next_2_2_sva);
  assign mux_77_nl = MUX_s_1_2_2(mux_76_nl, mux_69_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign mux_661_nl = MUX_s_1_2_2(or_tmp_87, or_dcpl_75, and_766_cse);
  assign mux_472_nl = MUX_s_1_2_2(mux_661_nl, or_dcpl_75, and_740_cse);
  assign mux_466_nl = MUX_s_1_2_2(mux_472_nl, or_dcpl_75, and_767_cse);
  assign mux_65_nl = MUX_s_1_2_2(mux_466_nl, or_dcpl_75, and_738_cse);
  assign mux_68_nl = MUX_s_1_2_2(mux_65_nl, or_dcpl_75, weight_mem_read_arbxbar_arbiters_next_2_6_sva);
  assign mux_78_nl = MUX_s_1_2_2(mux_77_nl, mux_68_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign mux_506_nl = MUX_s_1_2_2(or_tmp_87, or_dcpl_75, and_766_cse);
  assign mux_478_nl = MUX_s_1_2_2(mux_506_nl, or_dcpl_75, and_740_cse);
  assign mux_477_nl = MUX_s_1_2_2(mux_478_nl, or_dcpl_75, and_767_cse);
  assign mux_476_nl = MUX_s_1_2_2(mux_477_nl, or_dcpl_75, and_738_cse);
  assign mux_66_nl = MUX_s_1_2_2(mux_476_nl, or_dcpl_75, and_768_cse);
  assign mux_67_nl = MUX_s_1_2_2(mux_66_nl, or_dcpl_75, weight_mem_read_arbxbar_arbiters_next_2_1_sva);
  assign mux_79_nl = MUX_s_1_2_2(mux_78_nl, mux_67_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign or_256_nl = (~(and_769_cse | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1))
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_80_nl = MUX_s_1_2_2(mux_79_nl, or_256_nl, while_stage_0_5);
  assign nor_503_nl = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]));
  assign mux_86_nl = MUX_s_1_2_2(nor_503_nl, mux_tmp_84, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign and_267_nl = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) & mux_tmp_84;
  assign mux_85_nl = MUX_s_1_2_2(and_267_nl, nor_tmp_29, weight_mem_read_arbxbar_arbiters_next_1_1_sva);
  assign mux_87_nl = MUX_s_1_2_2(mux_86_nl, mux_85_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign mux_88_nl = MUX_s_1_2_2(mux_87_nl, nor_tmp_29, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign or_270_nl = (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | mux_88_nl;
  assign or_266_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(or_dcpl_40 | and_803_cse));
  assign mux_89_nl = MUX_s_1_2_2(or_270_nl, or_266_nl, while_stage_0_5);
  assign or_279_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_tmp
      | or_tmp_104;
  assign or_876_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_tmp
      | nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_5_mux_mx0w3))
      | or_tmp_104;
  assign nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_nl
      = MUX_s_1_2_2(operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_tmp);
  assign mux_91_nl = MUX_s_1_2_2(or_279_nl, or_876_nl, nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_nl);
  assign or_277_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp
      | or_tmp_104;
  assign nand_2_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp
      & (~ or_tmp_104));
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_1_nl
      = MUX_s_1_2_2(nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_3_mux_mx0w1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_mx0w0,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp);
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_37_nl
      = MUX_s_1_2_2(operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_tmp);
  assign nor_35_nl = ~(nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_1_nl
      | (~ nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_37_nl));
  assign mux_90_nl = MUX_s_1_2_2(or_277_nl, nand_2_nl, nor_35_nl);
  assign mux_92_nl = MUX_s_1_2_2(mux_91_nl, mux_90_nl, weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign or_274_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp
      | and_804_cse));
  assign mux_93_nl = MUX_s_1_2_2(mux_92_nl, or_274_nl, while_stage_0_5);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl
      = pe_manager_base_input_sva_mx1_7_0 & ({{7{and_319_cse}}, and_319_cse}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_1_nl
      = MUX_v_8_2_2(8'b00000000, pe_config_input_counter_sva_mx1, PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl
      = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]), pe_config_is_zero_first_sva_mx1,
      PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_27_nl
      = MUX_s_1_2_2(PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl,
      pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_or_5_cse_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_135_nl = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b110)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_142_nl = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_132_nl = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b011)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_1_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_1_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b101)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_1_tmp;
  assign mux_95_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, (~ pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign PECore_RunScale_if_for_1_scaled_val_mul_1_nl = (accum_vector_data_0_19_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_6_scaled_val_mul_1_nl = (accum_vector_data_5_19_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_7_scaled_val_mul_1_nl = (accum_vector_data_6_19_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_8_scaled_val_mul_1_nl = (accum_vector_data_7_19_0_sva)
      * 8'b10100111;
  assign act_port_reg_operator_for_act_port_reg_operator_for_and_nl = MUX_v_17_2_2(17'b00000000000000000,
      act_port_reg_data_16_0_sva_dfm_3, fsm_output);
  assign act_port_reg_operator_for_act_port_reg_operator_for_and_1_nl = MUX_v_17_2_2(17'b00000000000000000,
      act_port_reg_data_176_160_sva_dfm_3, fsm_output);
  assign act_port_reg_operator_for_act_port_reg_operator_for_and_2_nl = MUX_v_17_2_2(17'b00000000000000000,
      act_port_reg_data_208_192_sva_dfm_3, fsm_output);
  assign act_port_reg_operator_for_act_port_reg_operator_for_and_3_nl = MUX_v_17_2_2(17'b00000000000000000,
      act_port_reg_data_240_224_sva_dfm_3, fsm_output);
  assign nl_ProductSum_for_acc_40_itm_1  = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_29_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_28_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_27_z);
  assign nl_ProductSum_for_acc_41_itm_1  = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_26_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_25_z);
  assign nl_ProductSum_for_acc_24_itm_1  = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_61_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_60_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_59_z);
  assign nl_ProductSum_for_acc_25_itm_1  = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_58_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_57_z);
  assign nl_ProductSum_for_acc_50_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_8_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_7_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_6_z);
  assign ProductSum_for_acc_50_nl = nl_ProductSum_for_acc_50_nl[19:0];
  assign nl_ProductSum_for_acc_51_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_5_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_4_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_3_z);
  assign ProductSum_for_acc_51_nl = nl_ProductSum_for_acc_51_nl[19:0];
  assign nl_ProductSum_for_acc_52_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_2_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_1_z);
  assign ProductSum_for_acc_52_nl = nl_ProductSum_for_acc_52_nl[18:0];
  assign nl_ProductSum_for_acc_nl = ProductSum_for_acc_50_nl + ProductSum_for_acc_51_nl
      + conv_u2s_19_20(ProductSum_for_acc_52_nl);
  assign ProductSum_for_acc_nl = nl_ProductSum_for_acc_nl[19:0];
  assign PECore_UpdateFSM_switch_lp_not_37_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign nl_ProductSum_for_acc_47_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_16_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_15_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_14_z);
  assign ProductSum_for_acc_47_nl = nl_ProductSum_for_acc_47_nl[19:0];
  assign nl_ProductSum_for_acc_48_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_13_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_12_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_11_z);
  assign ProductSum_for_acc_48_nl = nl_ProductSum_for_acc_48_nl[19:0];
  assign nl_ProductSum_for_acc_49_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_10_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_9_z);
  assign ProductSum_for_acc_49_nl = nl_ProductSum_for_acc_49_nl[18:0];
  assign nl_ProductSum_for_acc_46_nl = ProductSum_for_acc_47_nl + ProductSum_for_acc_48_nl
      + conv_u2s_19_20(ProductSum_for_acc_49_nl);
  assign ProductSum_for_acc_46_nl = nl_ProductSum_for_acc_46_nl[19:0];
  assign PECore_UpdateFSM_switch_lp_not_23_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign nl_ProductSum_for_acc_43_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_24_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_23_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_22_z);
  assign ProductSum_for_acc_43_nl = nl_ProductSum_for_acc_43_nl[19:0];
  assign nl_ProductSum_for_acc_44_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_21_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_20_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_19_z);
  assign ProductSum_for_acc_44_nl = nl_ProductSum_for_acc_44_nl[19:0];
  assign nl_ProductSum_for_acc_45_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_18_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_17_z);
  assign ProductSum_for_acc_45_nl = nl_ProductSum_for_acc_45_nl[18:0];
  assign nl_ProductSum_for_acc_42_nl = ProductSum_for_acc_43_nl + ProductSum_for_acc_44_nl
      + conv_u2s_19_20(ProductSum_for_acc_45_nl);
  assign ProductSum_for_acc_42_nl = nl_ProductSum_for_acc_42_nl[19:0];
  assign PECore_UpdateFSM_switch_lp_not_38_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign nl_ProductSum_for_acc_35_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_40_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_39_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_38_z);
  assign ProductSum_for_acc_35_nl = nl_ProductSum_for_acc_35_nl[19:0];
  assign nl_ProductSum_for_acc_36_nl = conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_37_z)
      + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_36_z) + conv_u2u_18_20(Datapath_for_4_ProductSum_for_acc_9_cmp_35_z);
  assign ProductSum_for_acc_36_nl = nl_ProductSum_for_acc_36_nl[19:0];
  assign nl_ProductSum_for_acc_37_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_34_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_9_cmp_33_z);
  assign ProductSum_for_acc_37_nl = nl_ProductSum_for_acc_37_nl[18:0];
  assign nl_ProductSum_for_acc_34_nl = ProductSum_for_acc_35_nl + ProductSum_for_acc_36_nl
      + conv_u2s_19_20(ProductSum_for_acc_37_nl);
  assign ProductSum_for_acc_34_nl = nl_ProductSum_for_acc_34_nl[19:0];
  assign PECore_UpdateFSM_switch_lp_not_39_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign and_1206_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & fsm_output;
  assign input_mem_banks_read_1_for_mux_nl = MUX_v_8_2_2(input_read_addrs_sva_1_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4,
      and_1206_nl);
  assign and_693_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & weight_mem_run_3_for_land_5_lpi_1_dfm_2;
  assign nor_612_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign weight_port_read_out_data_mux_144_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_23_mx0w2,
      (weight_port_read_out_data_0_7_sva_dfm_mx0w2[7]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_703_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign nor_616_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_248_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[15:8]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_248_nl);
  assign while_if_while_if_and_2_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:0])
      & ({{14{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & ({{14{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
  assign or_465_nl = or_dcpl_151 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) |
      (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | or_dcpl_284;
  assign or_317_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]);
  assign mux_105_nl = MUX_s_1_2_2(and_dcpl_197, or_317_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_2);
  assign and_805_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & rva_in_reg_rw_sva_3;
  assign mux_108_nl = MUX_s_1_2_2(or_1106_cse, and_805_nl, weight_mem_run_3_for_weight_mem_run_3_for_and_6_tmp);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_103_itm_1
      & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_31_itm_1
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2,
      pe_manager_base_weight_sva_mx3_0, PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2,
      (pe_manager_base_weight_sva_mx2[8]), PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl =
      (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl = MUX_s_1_2_2(pe_config_is_valid_sva,
      pe_manager_zero_active_sva, and_319_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl = MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1,
      (pe_manager_num_input_sva[0]), and_319_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_6_nl = MUX_v_4_2_2(pe_config_num_manager_sva,
      (pe_manager_base_bias_sva[3:0]), and_319_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl = MUX_v_7_2_2((pe_config_num_output_sva[6:0]),
      (pe_manager_base_bias_sva[14:8]), and_319_cse);
  assign mux1h_nl = MUX1HOT_v_4_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_7_4,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1[7:4]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[31:28]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[31:28]),
      weight_port_read_out_data_0_3_sva_mx0_7_4, {and_1147_cse , and_1148_cse , and_1149_cse
      , and_1150_cse , and_1151_cse , and_1152_cse , nor_626_cse});
  assign not_2446_nl = ~ or_dcpl;
  assign mux1h_8_nl = MUX1HOT_v_4_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1_3_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1[3:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[27:24]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[27:24]),
      weight_port_read_out_data_0_3_sva_mx0_3_0, {and_1147_cse , and_1148_cse , and_1149_cse
      , and_1150_cse , and_1151_cse , and_1152_cse , nor_626_cse});
  assign not_2368_nl = ~ or_dcpl;
  assign mux1h_11_nl = MUX1HOT_v_7_7_2((rva_out_reg_data_55_48_sva_dfm_1_5[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[14:8]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[14:8]),
      weight_port_read_out_data_0_1_sva_mx0_6_0, {and_1147_cse , and_1148_cse , and_1149_cse
      , and_1150_cse , and_1151_cse , and_1152_cse , nor_626_cse});
  assign not_2449_nl = ~ or_dcpl;
  assign mux1h_9_nl = MUX1HOT_v_2_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7_4[1:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_5_0[5:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1[5:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1[5:4]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[21:20]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[21:20]),
      weight_port_read_out_data_0_2_sva_mx0_5_4, {and_1155_ssc , and_1156_cse , and_1157_cse
      , and_1158_cse , and_1159_cse , and_1160_cse , nor_627_cse});
  assign not_2448_nl = ~ or_dcpl_296;
  assign mux1h_2_nl = MUX1HOT_s_1_7_2((rva_out_reg_data_55_48_sva_dfm_1_5[7]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[15]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[15]),
      weight_port_read_out_data_0_1_sva_mx0_7, {and_1147_cse , and_1148_cse , and_1149_cse
      , and_1150_cse , and_1151_cse , and_1152_cse , nor_626_cse});
  assign mux1h_1_nl = MUX1HOT_s_1_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7_4[3]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_7_6[1]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[23]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[23]),
      weight_port_read_out_data_0_2_sva_mx0_7, {and_1155_ssc , and_1156_cse , and_1157_cse
      , and_1158_cse , and_1159_cse , and_1160_cse , nor_627_cse});
  assign mux1h_15_nl = MUX1HOT_s_1_7_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7_4[2]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_7_6[0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1[6]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[22]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[22]),
      weight_port_read_out_data_0_2_sva_mx0_6, {and_1155_ssc , and_1156_cse , and_1157_cse
      , and_1158_cse , and_1159_cse , and_1160_cse , nor_627_cse});
  assign mux1h_10_nl = MUX1HOT_v_4_7_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_3_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1_5_0[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1[3:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[19:16]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[19:16]),
      weight_port_read_out_data_0_2_sva_mx0_3_0, {and_1155_ssc , and_1156_cse , and_1157_cse
      , and_1158_cse , and_1159_cse , and_1160_cse , nor_627_cse});
  assign not_2370_nl = ~ or_dcpl_296;
  assign weight_mem_banks_load_store_for_else_mux1h_61_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[47]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[47]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[47]),
      {and_dcpl_659 , and_dcpl_661 , and_dcpl_662});
  assign weight_mem_banks_load_store_for_else_mux1h_86_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[46:40]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[46:40]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[46:40]),
      rva_out_reg_data_62_56_sva_dfm_1_4, {and_dcpl_659 , and_dcpl_661 , and_dcpl_662
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2357_nl = ~ or_dcpl_300;
  assign weight_mem_banks_load_store_for_else_mux1h_66_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[39]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[39]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[39]),
      {and_dcpl_659 , and_dcpl_661 , and_dcpl_662});
  assign weight_mem_banks_load_store_for_else_mux1h_87_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[38:32]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[38:32]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[38:32]),
      rva_out_reg_data_46_40_sva_dfm_1_4, {and_dcpl_659 , and_dcpl_661 , and_dcpl_662
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2359_nl = ~ or_dcpl_300;
  assign weight_mem_banks_load_store_for_else_mux1h_71_nl = MUX1HOT_v_4_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[31:28]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[31:28]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[31:28]),
      {and_dcpl_659 , and_dcpl_661 , and_dcpl_662});
  assign not_2360_nl = ~ or_dcpl_300;
  assign weight_mem_banks_load_store_for_else_mux1h_88_nl = MUX1HOT_v_4_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[27:24]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[27:24]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[27:24]),
      rva_out_reg_data_35_32_sva_dfm_1_4, {and_dcpl_659 , and_dcpl_661 , and_dcpl_662
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2361_nl = ~ or_dcpl_300;
  assign weight_mem_banks_load_store_for_else_mux1h_76_nl = MUX1HOT_v_2_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[23:22]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[23:22]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[23:22]),
      {and_dcpl_659 , and_dcpl_661 , and_dcpl_662});
  assign not_2362_nl = ~ or_dcpl_300;
  assign weight_mem_banks_load_store_for_else_mux1h_89_nl = MUX1HOT_v_6_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[21:16]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[21:16]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[21:16]),
      rva_out_reg_data_30_25_sva_dfm_2, {and_dcpl_659 , and_dcpl_661 , and_dcpl_662
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2363_nl = ~ or_dcpl_300;
  assign weight_mem_banks_load_store_for_else_mux1h_80_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[15]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[15]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[15]),
      {and_dcpl_659 , and_dcpl_661 , and_dcpl_662});
  assign weight_mem_banks_load_store_for_else_mux1h_90_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[14:8]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[14:8]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[14:8]),
      rva_out_reg_data_23_17_sva_dfm_2, {and_dcpl_659 , and_dcpl_661 , and_dcpl_662
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2365_nl = ~ or_dcpl_300;
  assign weight_mem_banks_load_store_for_else_mux1h_85_nl = MUX1HOT_s_1_5_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[7]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[7]), (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[7]),
      (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[7]), (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[7]),
      {and_677_ssc , and_678_ssc , and_680_ssc , and_683_ssc , and_686_ssc});
  assign weight_mem_banks_load_store_for_else_or_nl = weight_mem_banks_load_store_for_else_mux1h_85_nl
      | and_676_ssc;
  assign mux_493_nl = MUX_s_1_2_2(weight_mem_banks_load_store_for_else_or_nl, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[7]),
      or_dcpl_301);
  assign and_687_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign weight_mem_banks_load_store_for_else_mux1h_91_nl = MUX1HOT_v_7_6_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[6:0]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[6:0]), (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[6:0]),
      (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[6:0]), (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[6:0]),
      rva_out_reg_data_15_9_sva_dfm_4, {and_677_ssc , and_678_ssc , and_680_ssc ,
      and_683_ssc , and_686_ssc , and_687_nl});
  assign weight_mem_banks_load_store_for_else_or_1_nl = MUX_v_7_2_2(weight_mem_banks_load_store_for_else_mux1h_91_nl,
      7'b1111111, and_676_ssc);
  assign mux_494_nl = MUX_v_7_2_2(weight_mem_banks_load_store_for_else_or_1_nl, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[6:0]),
      or_dcpl_301);
  assign not_2367_nl = ~ and_dcpl_737;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[103:100]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_268_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_237_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_130_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[99:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_237_nl);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_nl
      = (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[95]) & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]));
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_128_nl
      = (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[94]) & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]));
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_265_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_135_nl
      = MUX_v_2_2_2(2'b00, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[93:92]), weight_mem_write_arbxbar_xbar_for_1_for_not_265_nl);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_nl
      = (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[87]) & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]));
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_136_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[91:88]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_266_nl);
  assign nor_745_nl = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_2 | (~ mux_tmp_560));
  assign mux_605_nl = MUX_s_1_2_2(mux_tmp_560, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_606_nl = MUX_s_1_2_2(nor_745_nl, mux_605_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_607_nl = MUX_s_1_2_2(mux_tmp_560, mux_606_nl, while_stage_0_6);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_267_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_129_nl
      = MUX_v_7_2_2(7'b0000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[86:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_267_nl);
  assign nor_746_nl = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_2 | (~ mux_tmp_567));
  assign mux_612_nl = MUX_s_1_2_2(mux_tmp_567, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_613_nl = MUX_s_1_2_2(nor_746_nl, mux_612_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_614_nl = MUX_s_1_2_2(mux_tmp_567, mux_613_nl, while_stage_0_6);
  assign or_1188_nl = reg_weight_mem_run_3_for_5_and_152_itm_2_cse | reg_weight_mem_run_3_for_5_and_151_itm_2_cse
      | weight_mem_run_3_for_5_and_150_itm_2 | reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      | weight_mem_run_3_for_5_and_148_itm_2 | reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_146_itm_2_cse | weight_mem_run_3_for_5_and_145_cse;
  assign or_1185_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2;
  assign or_1184_nl = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2;
  assign mux_615_nl = MUX_s_1_2_2(or_1185_nl, or_1184_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign or_1183_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_33_itm_2;
  assign mux_616_nl = MUX_s_1_2_2(mux_615_nl, or_1183_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_1186_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_239_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 | (crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & mux_616_nl);
  assign mux_617_nl = MUX_s_1_2_2(or_1188_nl, or_1186_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_nl
      = (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[119]) & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]));
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_nl
      = (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[111]) & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]));

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_9_2;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [8:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_8_2;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [7:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    result = result | (input_5 & {11{sel[5]}});
    result = result | (input_6 & {11{sel[6]}});
    result = result | (input_7 & {11{sel[7]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function automatic [127:0] MUX1HOT_v_128_3_2;
    input [127:0] input_2;
    input [127:0] input_1;
    input [127:0] input_0;
    input [2:0] sel;
    reg [127:0] result;
  begin
    result = input_0 & {128{sel[0]}};
    result = result | (input_1 & {128{sel[1]}});
    result = result | (input_2 & {128{sel[2]}});
    MUX1HOT_v_128_3_2 = result;
  end
  endfunction


  function automatic [16:0] MUX1HOT_v_17_3_2;
    input [16:0] input_2;
    input [16:0] input_1;
    input [16:0] input_0;
    input [2:0] sel;
    reg [16:0] result;
  begin
    result = input_0 & {17{sel[0]}};
    result = result | (input_1 & {17{sel[1]}});
    result = result | (input_2 & {17{sel[2]}});
    MUX1HOT_v_17_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_7_2;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [6:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    MUX1HOT_v_2_7_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_7_2;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [6:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    MUX1HOT_v_4_7_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_6_2;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [5:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    MUX1HOT_v_7_6_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_7_2;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [6:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    result = result | (input_6 & {7{sel[6]}});
    MUX1HOT_v_7_7_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_9_2;
    input [6:0] input_8;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [8:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    result = result | (input_6 & {7{sel[6]}});
    result = result | (input_7 & {7{sel[7]}});
    result = result | (input_8 & {7{sel[8]}});
    MUX1HOT_v_7_9_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_7_2;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [6:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    MUX1HOT_v_8_7_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_8_2;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [7:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    MUX1HOT_v_8_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_9_2;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [8:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    result = result | (input_8 & {8{sel[8]}});
    MUX1HOT_v_8_9_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_8_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input [2:0] sel;
    reg  result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_s_1_8_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_8_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [10:0] input_2;
    input [10:0] input_3;
    input [10:0] input_4;
    input [10:0] input_5;
    input [10:0] input_6;
    input [10:0] input_7;
    input [2:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_11_8_2 = result;
  end
  endfunction


  function automatic [119:0] MUX_v_120_2_2;
    input [119:0] input_0;
    input [119:0] input_1;
    input  sel;
    reg [119:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_120_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_256_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [127:0] input_2;
    input [127:0] input_3;
    input [127:0] input_4;
    input [127:0] input_5;
    input [127:0] input_6;
    input [127:0] input_7;
    input [127:0] input_8;
    input [127:0] input_9;
    input [127:0] input_10;
    input [127:0] input_11;
    input [127:0] input_12;
    input [127:0] input_13;
    input [127:0] input_14;
    input [127:0] input_15;
    input [127:0] input_16;
    input [127:0] input_17;
    input [127:0] input_18;
    input [127:0] input_19;
    input [127:0] input_20;
    input [127:0] input_21;
    input [127:0] input_22;
    input [127:0] input_23;
    input [127:0] input_24;
    input [127:0] input_25;
    input [127:0] input_26;
    input [127:0] input_27;
    input [127:0] input_28;
    input [127:0] input_29;
    input [127:0] input_30;
    input [127:0] input_31;
    input [127:0] input_32;
    input [127:0] input_33;
    input [127:0] input_34;
    input [127:0] input_35;
    input [127:0] input_36;
    input [127:0] input_37;
    input [127:0] input_38;
    input [127:0] input_39;
    input [127:0] input_40;
    input [127:0] input_41;
    input [127:0] input_42;
    input [127:0] input_43;
    input [127:0] input_44;
    input [127:0] input_45;
    input [127:0] input_46;
    input [127:0] input_47;
    input [127:0] input_48;
    input [127:0] input_49;
    input [127:0] input_50;
    input [127:0] input_51;
    input [127:0] input_52;
    input [127:0] input_53;
    input [127:0] input_54;
    input [127:0] input_55;
    input [127:0] input_56;
    input [127:0] input_57;
    input [127:0] input_58;
    input [127:0] input_59;
    input [127:0] input_60;
    input [127:0] input_61;
    input [127:0] input_62;
    input [127:0] input_63;
    input [127:0] input_64;
    input [127:0] input_65;
    input [127:0] input_66;
    input [127:0] input_67;
    input [127:0] input_68;
    input [127:0] input_69;
    input [127:0] input_70;
    input [127:0] input_71;
    input [127:0] input_72;
    input [127:0] input_73;
    input [127:0] input_74;
    input [127:0] input_75;
    input [127:0] input_76;
    input [127:0] input_77;
    input [127:0] input_78;
    input [127:0] input_79;
    input [127:0] input_80;
    input [127:0] input_81;
    input [127:0] input_82;
    input [127:0] input_83;
    input [127:0] input_84;
    input [127:0] input_85;
    input [127:0] input_86;
    input [127:0] input_87;
    input [127:0] input_88;
    input [127:0] input_89;
    input [127:0] input_90;
    input [127:0] input_91;
    input [127:0] input_92;
    input [127:0] input_93;
    input [127:0] input_94;
    input [127:0] input_95;
    input [127:0] input_96;
    input [127:0] input_97;
    input [127:0] input_98;
    input [127:0] input_99;
    input [127:0] input_100;
    input [127:0] input_101;
    input [127:0] input_102;
    input [127:0] input_103;
    input [127:0] input_104;
    input [127:0] input_105;
    input [127:0] input_106;
    input [127:0] input_107;
    input [127:0] input_108;
    input [127:0] input_109;
    input [127:0] input_110;
    input [127:0] input_111;
    input [127:0] input_112;
    input [127:0] input_113;
    input [127:0] input_114;
    input [127:0] input_115;
    input [127:0] input_116;
    input [127:0] input_117;
    input [127:0] input_118;
    input [127:0] input_119;
    input [127:0] input_120;
    input [127:0] input_121;
    input [127:0] input_122;
    input [127:0] input_123;
    input [127:0] input_124;
    input [127:0] input_125;
    input [127:0] input_126;
    input [127:0] input_127;
    input [127:0] input_128;
    input [127:0] input_129;
    input [127:0] input_130;
    input [127:0] input_131;
    input [127:0] input_132;
    input [127:0] input_133;
    input [127:0] input_134;
    input [127:0] input_135;
    input [127:0] input_136;
    input [127:0] input_137;
    input [127:0] input_138;
    input [127:0] input_139;
    input [127:0] input_140;
    input [127:0] input_141;
    input [127:0] input_142;
    input [127:0] input_143;
    input [127:0] input_144;
    input [127:0] input_145;
    input [127:0] input_146;
    input [127:0] input_147;
    input [127:0] input_148;
    input [127:0] input_149;
    input [127:0] input_150;
    input [127:0] input_151;
    input [127:0] input_152;
    input [127:0] input_153;
    input [127:0] input_154;
    input [127:0] input_155;
    input [127:0] input_156;
    input [127:0] input_157;
    input [127:0] input_158;
    input [127:0] input_159;
    input [127:0] input_160;
    input [127:0] input_161;
    input [127:0] input_162;
    input [127:0] input_163;
    input [127:0] input_164;
    input [127:0] input_165;
    input [127:0] input_166;
    input [127:0] input_167;
    input [127:0] input_168;
    input [127:0] input_169;
    input [127:0] input_170;
    input [127:0] input_171;
    input [127:0] input_172;
    input [127:0] input_173;
    input [127:0] input_174;
    input [127:0] input_175;
    input [127:0] input_176;
    input [127:0] input_177;
    input [127:0] input_178;
    input [127:0] input_179;
    input [127:0] input_180;
    input [127:0] input_181;
    input [127:0] input_182;
    input [127:0] input_183;
    input [127:0] input_184;
    input [127:0] input_185;
    input [127:0] input_186;
    input [127:0] input_187;
    input [127:0] input_188;
    input [127:0] input_189;
    input [127:0] input_190;
    input [127:0] input_191;
    input [127:0] input_192;
    input [127:0] input_193;
    input [127:0] input_194;
    input [127:0] input_195;
    input [127:0] input_196;
    input [127:0] input_197;
    input [127:0] input_198;
    input [127:0] input_199;
    input [127:0] input_200;
    input [127:0] input_201;
    input [127:0] input_202;
    input [127:0] input_203;
    input [127:0] input_204;
    input [127:0] input_205;
    input [127:0] input_206;
    input [127:0] input_207;
    input [127:0] input_208;
    input [127:0] input_209;
    input [127:0] input_210;
    input [127:0] input_211;
    input [127:0] input_212;
    input [127:0] input_213;
    input [127:0] input_214;
    input [127:0] input_215;
    input [127:0] input_216;
    input [127:0] input_217;
    input [127:0] input_218;
    input [127:0] input_219;
    input [127:0] input_220;
    input [127:0] input_221;
    input [127:0] input_222;
    input [127:0] input_223;
    input [127:0] input_224;
    input [127:0] input_225;
    input [127:0] input_226;
    input [127:0] input_227;
    input [127:0] input_228;
    input [127:0] input_229;
    input [127:0] input_230;
    input [127:0] input_231;
    input [127:0] input_232;
    input [127:0] input_233;
    input [127:0] input_234;
    input [127:0] input_235;
    input [127:0] input_236;
    input [127:0] input_237;
    input [127:0] input_238;
    input [127:0] input_239;
    input [127:0] input_240;
    input [127:0] input_241;
    input [127:0] input_242;
    input [127:0] input_243;
    input [127:0] input_244;
    input [127:0] input_245;
    input [127:0] input_246;
    input [127:0] input_247;
    input [127:0] input_248;
    input [127:0] input_249;
    input [127:0] input_250;
    input [127:0] input_251;
    input [127:0] input_252;
    input [127:0] input_253;
    input [127:0] input_254;
    input [127:0] input_255;
    input [7:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      8'b00000000 : begin
        result = input_0;
      end
      8'b00000001 : begin
        result = input_1;
      end
      8'b00000010 : begin
        result = input_2;
      end
      8'b00000011 : begin
        result = input_3;
      end
      8'b00000100 : begin
        result = input_4;
      end
      8'b00000101 : begin
        result = input_5;
      end
      8'b00000110 : begin
        result = input_6;
      end
      8'b00000111 : begin
        result = input_7;
      end
      8'b00001000 : begin
        result = input_8;
      end
      8'b00001001 : begin
        result = input_9;
      end
      8'b00001010 : begin
        result = input_10;
      end
      8'b00001011 : begin
        result = input_11;
      end
      8'b00001100 : begin
        result = input_12;
      end
      8'b00001101 : begin
        result = input_13;
      end
      8'b00001110 : begin
        result = input_14;
      end
      8'b00001111 : begin
        result = input_15;
      end
      8'b00010000 : begin
        result = input_16;
      end
      8'b00010001 : begin
        result = input_17;
      end
      8'b00010010 : begin
        result = input_18;
      end
      8'b00010011 : begin
        result = input_19;
      end
      8'b00010100 : begin
        result = input_20;
      end
      8'b00010101 : begin
        result = input_21;
      end
      8'b00010110 : begin
        result = input_22;
      end
      8'b00010111 : begin
        result = input_23;
      end
      8'b00011000 : begin
        result = input_24;
      end
      8'b00011001 : begin
        result = input_25;
      end
      8'b00011010 : begin
        result = input_26;
      end
      8'b00011011 : begin
        result = input_27;
      end
      8'b00011100 : begin
        result = input_28;
      end
      8'b00011101 : begin
        result = input_29;
      end
      8'b00011110 : begin
        result = input_30;
      end
      8'b00011111 : begin
        result = input_31;
      end
      8'b00100000 : begin
        result = input_32;
      end
      8'b00100001 : begin
        result = input_33;
      end
      8'b00100010 : begin
        result = input_34;
      end
      8'b00100011 : begin
        result = input_35;
      end
      8'b00100100 : begin
        result = input_36;
      end
      8'b00100101 : begin
        result = input_37;
      end
      8'b00100110 : begin
        result = input_38;
      end
      8'b00100111 : begin
        result = input_39;
      end
      8'b00101000 : begin
        result = input_40;
      end
      8'b00101001 : begin
        result = input_41;
      end
      8'b00101010 : begin
        result = input_42;
      end
      8'b00101011 : begin
        result = input_43;
      end
      8'b00101100 : begin
        result = input_44;
      end
      8'b00101101 : begin
        result = input_45;
      end
      8'b00101110 : begin
        result = input_46;
      end
      8'b00101111 : begin
        result = input_47;
      end
      8'b00110000 : begin
        result = input_48;
      end
      8'b00110001 : begin
        result = input_49;
      end
      8'b00110010 : begin
        result = input_50;
      end
      8'b00110011 : begin
        result = input_51;
      end
      8'b00110100 : begin
        result = input_52;
      end
      8'b00110101 : begin
        result = input_53;
      end
      8'b00110110 : begin
        result = input_54;
      end
      8'b00110111 : begin
        result = input_55;
      end
      8'b00111000 : begin
        result = input_56;
      end
      8'b00111001 : begin
        result = input_57;
      end
      8'b00111010 : begin
        result = input_58;
      end
      8'b00111011 : begin
        result = input_59;
      end
      8'b00111100 : begin
        result = input_60;
      end
      8'b00111101 : begin
        result = input_61;
      end
      8'b00111110 : begin
        result = input_62;
      end
      8'b00111111 : begin
        result = input_63;
      end
      8'b01000000 : begin
        result = input_64;
      end
      8'b01000001 : begin
        result = input_65;
      end
      8'b01000010 : begin
        result = input_66;
      end
      8'b01000011 : begin
        result = input_67;
      end
      8'b01000100 : begin
        result = input_68;
      end
      8'b01000101 : begin
        result = input_69;
      end
      8'b01000110 : begin
        result = input_70;
      end
      8'b01000111 : begin
        result = input_71;
      end
      8'b01001000 : begin
        result = input_72;
      end
      8'b01001001 : begin
        result = input_73;
      end
      8'b01001010 : begin
        result = input_74;
      end
      8'b01001011 : begin
        result = input_75;
      end
      8'b01001100 : begin
        result = input_76;
      end
      8'b01001101 : begin
        result = input_77;
      end
      8'b01001110 : begin
        result = input_78;
      end
      8'b01001111 : begin
        result = input_79;
      end
      8'b01010000 : begin
        result = input_80;
      end
      8'b01010001 : begin
        result = input_81;
      end
      8'b01010010 : begin
        result = input_82;
      end
      8'b01010011 : begin
        result = input_83;
      end
      8'b01010100 : begin
        result = input_84;
      end
      8'b01010101 : begin
        result = input_85;
      end
      8'b01010110 : begin
        result = input_86;
      end
      8'b01010111 : begin
        result = input_87;
      end
      8'b01011000 : begin
        result = input_88;
      end
      8'b01011001 : begin
        result = input_89;
      end
      8'b01011010 : begin
        result = input_90;
      end
      8'b01011011 : begin
        result = input_91;
      end
      8'b01011100 : begin
        result = input_92;
      end
      8'b01011101 : begin
        result = input_93;
      end
      8'b01011110 : begin
        result = input_94;
      end
      8'b01011111 : begin
        result = input_95;
      end
      8'b01100000 : begin
        result = input_96;
      end
      8'b01100001 : begin
        result = input_97;
      end
      8'b01100010 : begin
        result = input_98;
      end
      8'b01100011 : begin
        result = input_99;
      end
      8'b01100100 : begin
        result = input_100;
      end
      8'b01100101 : begin
        result = input_101;
      end
      8'b01100110 : begin
        result = input_102;
      end
      8'b01100111 : begin
        result = input_103;
      end
      8'b01101000 : begin
        result = input_104;
      end
      8'b01101001 : begin
        result = input_105;
      end
      8'b01101010 : begin
        result = input_106;
      end
      8'b01101011 : begin
        result = input_107;
      end
      8'b01101100 : begin
        result = input_108;
      end
      8'b01101101 : begin
        result = input_109;
      end
      8'b01101110 : begin
        result = input_110;
      end
      8'b01101111 : begin
        result = input_111;
      end
      8'b01110000 : begin
        result = input_112;
      end
      8'b01110001 : begin
        result = input_113;
      end
      8'b01110010 : begin
        result = input_114;
      end
      8'b01110011 : begin
        result = input_115;
      end
      8'b01110100 : begin
        result = input_116;
      end
      8'b01110101 : begin
        result = input_117;
      end
      8'b01110110 : begin
        result = input_118;
      end
      8'b01110111 : begin
        result = input_119;
      end
      8'b01111000 : begin
        result = input_120;
      end
      8'b01111001 : begin
        result = input_121;
      end
      8'b01111010 : begin
        result = input_122;
      end
      8'b01111011 : begin
        result = input_123;
      end
      8'b01111100 : begin
        result = input_124;
      end
      8'b01111101 : begin
        result = input_125;
      end
      8'b01111110 : begin
        result = input_126;
      end
      8'b01111111 : begin
        result = input_127;
      end
      8'b10000000 : begin
        result = input_128;
      end
      8'b10000001 : begin
        result = input_129;
      end
      8'b10000010 : begin
        result = input_130;
      end
      8'b10000011 : begin
        result = input_131;
      end
      8'b10000100 : begin
        result = input_132;
      end
      8'b10000101 : begin
        result = input_133;
      end
      8'b10000110 : begin
        result = input_134;
      end
      8'b10000111 : begin
        result = input_135;
      end
      8'b10001000 : begin
        result = input_136;
      end
      8'b10001001 : begin
        result = input_137;
      end
      8'b10001010 : begin
        result = input_138;
      end
      8'b10001011 : begin
        result = input_139;
      end
      8'b10001100 : begin
        result = input_140;
      end
      8'b10001101 : begin
        result = input_141;
      end
      8'b10001110 : begin
        result = input_142;
      end
      8'b10001111 : begin
        result = input_143;
      end
      8'b10010000 : begin
        result = input_144;
      end
      8'b10010001 : begin
        result = input_145;
      end
      8'b10010010 : begin
        result = input_146;
      end
      8'b10010011 : begin
        result = input_147;
      end
      8'b10010100 : begin
        result = input_148;
      end
      8'b10010101 : begin
        result = input_149;
      end
      8'b10010110 : begin
        result = input_150;
      end
      8'b10010111 : begin
        result = input_151;
      end
      8'b10011000 : begin
        result = input_152;
      end
      8'b10011001 : begin
        result = input_153;
      end
      8'b10011010 : begin
        result = input_154;
      end
      8'b10011011 : begin
        result = input_155;
      end
      8'b10011100 : begin
        result = input_156;
      end
      8'b10011101 : begin
        result = input_157;
      end
      8'b10011110 : begin
        result = input_158;
      end
      8'b10011111 : begin
        result = input_159;
      end
      8'b10100000 : begin
        result = input_160;
      end
      8'b10100001 : begin
        result = input_161;
      end
      8'b10100010 : begin
        result = input_162;
      end
      8'b10100011 : begin
        result = input_163;
      end
      8'b10100100 : begin
        result = input_164;
      end
      8'b10100101 : begin
        result = input_165;
      end
      8'b10100110 : begin
        result = input_166;
      end
      8'b10100111 : begin
        result = input_167;
      end
      8'b10101000 : begin
        result = input_168;
      end
      8'b10101001 : begin
        result = input_169;
      end
      8'b10101010 : begin
        result = input_170;
      end
      8'b10101011 : begin
        result = input_171;
      end
      8'b10101100 : begin
        result = input_172;
      end
      8'b10101101 : begin
        result = input_173;
      end
      8'b10101110 : begin
        result = input_174;
      end
      8'b10101111 : begin
        result = input_175;
      end
      8'b10110000 : begin
        result = input_176;
      end
      8'b10110001 : begin
        result = input_177;
      end
      8'b10110010 : begin
        result = input_178;
      end
      8'b10110011 : begin
        result = input_179;
      end
      8'b10110100 : begin
        result = input_180;
      end
      8'b10110101 : begin
        result = input_181;
      end
      8'b10110110 : begin
        result = input_182;
      end
      8'b10110111 : begin
        result = input_183;
      end
      8'b10111000 : begin
        result = input_184;
      end
      8'b10111001 : begin
        result = input_185;
      end
      8'b10111010 : begin
        result = input_186;
      end
      8'b10111011 : begin
        result = input_187;
      end
      8'b10111100 : begin
        result = input_188;
      end
      8'b10111101 : begin
        result = input_189;
      end
      8'b10111110 : begin
        result = input_190;
      end
      8'b10111111 : begin
        result = input_191;
      end
      8'b11000000 : begin
        result = input_192;
      end
      8'b11000001 : begin
        result = input_193;
      end
      8'b11000010 : begin
        result = input_194;
      end
      8'b11000011 : begin
        result = input_195;
      end
      8'b11000100 : begin
        result = input_196;
      end
      8'b11000101 : begin
        result = input_197;
      end
      8'b11000110 : begin
        result = input_198;
      end
      8'b11000111 : begin
        result = input_199;
      end
      8'b11001000 : begin
        result = input_200;
      end
      8'b11001001 : begin
        result = input_201;
      end
      8'b11001010 : begin
        result = input_202;
      end
      8'b11001011 : begin
        result = input_203;
      end
      8'b11001100 : begin
        result = input_204;
      end
      8'b11001101 : begin
        result = input_205;
      end
      8'b11001110 : begin
        result = input_206;
      end
      8'b11001111 : begin
        result = input_207;
      end
      8'b11010000 : begin
        result = input_208;
      end
      8'b11010001 : begin
        result = input_209;
      end
      8'b11010010 : begin
        result = input_210;
      end
      8'b11010011 : begin
        result = input_211;
      end
      8'b11010100 : begin
        result = input_212;
      end
      8'b11010101 : begin
        result = input_213;
      end
      8'b11010110 : begin
        result = input_214;
      end
      8'b11010111 : begin
        result = input_215;
      end
      8'b11011000 : begin
        result = input_216;
      end
      8'b11011001 : begin
        result = input_217;
      end
      8'b11011010 : begin
        result = input_218;
      end
      8'b11011011 : begin
        result = input_219;
      end
      8'b11011100 : begin
        result = input_220;
      end
      8'b11011101 : begin
        result = input_221;
      end
      8'b11011110 : begin
        result = input_222;
      end
      8'b11011111 : begin
        result = input_223;
      end
      8'b11100000 : begin
        result = input_224;
      end
      8'b11100001 : begin
        result = input_225;
      end
      8'b11100010 : begin
        result = input_226;
      end
      8'b11100011 : begin
        result = input_227;
      end
      8'b11100100 : begin
        result = input_228;
      end
      8'b11100101 : begin
        result = input_229;
      end
      8'b11100110 : begin
        result = input_230;
      end
      8'b11100111 : begin
        result = input_231;
      end
      8'b11101000 : begin
        result = input_232;
      end
      8'b11101001 : begin
        result = input_233;
      end
      8'b11101010 : begin
        result = input_234;
      end
      8'b11101011 : begin
        result = input_235;
      end
      8'b11101100 : begin
        result = input_236;
      end
      8'b11101101 : begin
        result = input_237;
      end
      8'b11101110 : begin
        result = input_238;
      end
      8'b11101111 : begin
        result = input_239;
      end
      8'b11110000 : begin
        result = input_240;
      end
      8'b11110001 : begin
        result = input_241;
      end
      8'b11110010 : begin
        result = input_242;
      end
      8'b11110011 : begin
        result = input_243;
      end
      8'b11110100 : begin
        result = input_244;
      end
      8'b11110101 : begin
        result = input_245;
      end
      8'b11110110 : begin
        result = input_246;
      end
      8'b11110111 : begin
        result = input_247;
      end
      8'b11111000 : begin
        result = input_248;
      end
      8'b11111001 : begin
        result = input_249;
      end
      8'b11111010 : begin
        result = input_250;
      end
      8'b11111011 : begin
        result = input_251;
      end
      8'b11111100 : begin
        result = input_252;
      end
      8'b11111101 : begin
        result = input_253;
      end
      8'b11111110 : begin
        result = input_254;
      end
      default : begin
        result = input_255;
      end
    endcase
    MUX_v_128_256_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input  sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input  sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input  sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_8_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [1:0] input_2;
    input [1:0] input_3;
    input [1:0] input_4;
    input [1:0] input_5;
    input [1:0] input_6;
    input [1:0] input_7;
    input [2:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_2_8_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_8_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [2:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_4_8_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_8_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [6:0] input_2;
    input [6:0] input_3;
    input [6:0] input_4;
    input [6:0] input_5;
    input [6:0] input_6;
    input [6:0] input_7;
    input [2:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_7_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [16:0] readslicef_28_17_11;
    input [27:0] vector;
    reg [27:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_28_17_11 = tmp[16:0];
  end
  endfunction


  function automatic [10:0] signext_11_1;
    input  vector;
  begin
    signext_11_1= {{10{vector}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input  vector;
  begin
    signext_4_1= {{3{vector}}, vector};
  end
  endfunction


  function automatic [5:0] signext_6_1;
    input  vector;
  begin
    signext_6_1= {{5{vector}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input  vector;
  begin
    signext_7_1= {{6{vector}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [19:0] conv_u2s_19_20 ;
    input [18:0]  vector ;
  begin
    conv_u2s_19_20 =  {1'b0, vector};
  end
  endfunction


  function automatic [18:0] conv_u2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_u2u_18_19 = {1'b0, vector};
  end
  endfunction


  function automatic [19:0] conv_u2u_18_20 ;
    input [17:0]  vector ;
  begin
    conv_u2u_18_20 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore
// ------------------------------------------------------------------


module PECore (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [137:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_c;
  wire Datapath_for_4_ProductSum_for_acc_9_cmp_en;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_c;
  wire Datapath_for_4_ProductSum_for_acc_9_cmp_1_en;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_z;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_1 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_1_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_1_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_1_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_2 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_2_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_2_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_2_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_3 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_3_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_3_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_3_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_4 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_4_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_4_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_4_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_5 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_5_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_5_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_5_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_6 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_6_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_6_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_6_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_7 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_7_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_7_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_7_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_8 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_8_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_8_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_8_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_9 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_9_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_9_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_9_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_10 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_10_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_10_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_10_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_11 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_11_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_11_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_11_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_12 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_12_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_12_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_12_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_13 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_13_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_13_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_13_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_14 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_14_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_14_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_14_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_15 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_15_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_15_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_15_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_16 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_16_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_16_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_16_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_17 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_17_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_17_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_17_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_18 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_18_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_18_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_18_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_19 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_19_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_19_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_19_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_20 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_20_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_20_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_20_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_21 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_21_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_21_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_21_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_22 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_22_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_22_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_22_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_23 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_23_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_23_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_23_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_24 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_24_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_24_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_24_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_25 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_25_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_25_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_25_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_26 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_26_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_26_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_26_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_27 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_27_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_27_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_27_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_28 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_28_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_28_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_28_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_29 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_29_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_29_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_29_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_30 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_30_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_30_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_30_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_31 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_31_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_31_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_31_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_32 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_32_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_32_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_32_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_33 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_33_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_33_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_33_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_34 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_34_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_34_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_34_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_35 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_35_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_35_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_35_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_36 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_36_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_36_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_36_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_37 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_37_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_37_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_37_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_38 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_38_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_38_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_38_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_39 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_39_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_39_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_39_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_40 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_40_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_40_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_40_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_41 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_41_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_41_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_41_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_41_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_41_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_42 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_42_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_42_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_42_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_42_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_42_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_43 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_43_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_43_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_43_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_43_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_43_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_44 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_44_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_44_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_44_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_44_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_44_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_45 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_45_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_45_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_45_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_45_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_45_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_46 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_46_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_46_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_46_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_46_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_46_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_47 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_47_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_47_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_47_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_47_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_47_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_48 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_48_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_48_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_48_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_49 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_49_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_41_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_49_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_41_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_49_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_50 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_50_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_42_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_50_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_42_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_50_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_51 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_51_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_43_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_51_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_43_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_51_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_52 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_52_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_44_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_52_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_44_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_52_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_53 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_53_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_45_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_53_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_45_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_53_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_54 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_54_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_46_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_54_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_46_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_54_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_55 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_55_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_47_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_55_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_47_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_55_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_56 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_56_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_56_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_56_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_57 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_57_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_57_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_57_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_58 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_58_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_58_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_58_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_59 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_59_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_59_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_59_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_60 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_60_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_60_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_60_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_61 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_61_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_61_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_61_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_62 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_62_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_62_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_62_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_63 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_63_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_63_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_63_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_PECoreRun PECore_PECoreRun_inst (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_a(Datapath_for_4_ProductSum_for_acc_9_cmp_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_c(Datapath_for_4_ProductSum_for_acc_9_cmp_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_z(Datapath_for_4_ProductSum_for_acc_9_cmp_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_a(Datapath_for_4_ProductSum_for_acc_9_cmp_1_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_c(Datapath_for_4_ProductSum_for_acc_9_cmp_1_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_z(Datapath_for_4_ProductSum_for_acc_9_cmp_1_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_a(Datapath_for_4_ProductSum_for_acc_9_cmp_2_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_c(Datapath_for_4_ProductSum_for_acc_9_cmp_2_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_z(Datapath_for_4_ProductSum_for_acc_9_cmp_2_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_a(Datapath_for_4_ProductSum_for_acc_9_cmp_3_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_c(Datapath_for_4_ProductSum_for_acc_9_cmp_3_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_z(Datapath_for_4_ProductSum_for_acc_9_cmp_3_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_a(Datapath_for_4_ProductSum_for_acc_9_cmp_4_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_c(Datapath_for_4_ProductSum_for_acc_9_cmp_4_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_z(Datapath_for_4_ProductSum_for_acc_9_cmp_4_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_a(Datapath_for_4_ProductSum_for_acc_9_cmp_5_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_c(Datapath_for_4_ProductSum_for_acc_9_cmp_5_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_z(Datapath_for_4_ProductSum_for_acc_9_cmp_5_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_a(Datapath_for_4_ProductSum_for_acc_9_cmp_6_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_c(Datapath_for_4_ProductSum_for_acc_9_cmp_6_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_z(Datapath_for_4_ProductSum_for_acc_9_cmp_6_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_a(Datapath_for_4_ProductSum_for_acc_9_cmp_7_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_c(Datapath_for_4_ProductSum_for_acc_9_cmp_7_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_z(Datapath_for_4_ProductSum_for_acc_9_cmp_7_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_a(Datapath_for_4_ProductSum_for_acc_9_cmp_8_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_c(Datapath_for_4_ProductSum_for_acc_9_cmp_8_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_z(Datapath_for_4_ProductSum_for_acc_9_cmp_8_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_9_a(Datapath_for_4_ProductSum_for_acc_9_cmp_9_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_9_c(Datapath_for_4_ProductSum_for_acc_9_cmp_9_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_9_z(Datapath_for_4_ProductSum_for_acc_9_cmp_9_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_10_a(Datapath_for_4_ProductSum_for_acc_9_cmp_10_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_10_c(Datapath_for_4_ProductSum_for_acc_9_cmp_10_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_10_z(Datapath_for_4_ProductSum_for_acc_9_cmp_10_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_11_a(Datapath_for_4_ProductSum_for_acc_9_cmp_11_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_11_c(Datapath_for_4_ProductSum_for_acc_9_cmp_11_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_11_z(Datapath_for_4_ProductSum_for_acc_9_cmp_11_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_12_a(Datapath_for_4_ProductSum_for_acc_9_cmp_12_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_12_c(Datapath_for_4_ProductSum_for_acc_9_cmp_12_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_12_z(Datapath_for_4_ProductSum_for_acc_9_cmp_12_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_13_a(Datapath_for_4_ProductSum_for_acc_9_cmp_13_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_13_c(Datapath_for_4_ProductSum_for_acc_9_cmp_13_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_13_z(Datapath_for_4_ProductSum_for_acc_9_cmp_13_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_14_a(Datapath_for_4_ProductSum_for_acc_9_cmp_14_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_14_c(Datapath_for_4_ProductSum_for_acc_9_cmp_14_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_14_z(Datapath_for_4_ProductSum_for_acc_9_cmp_14_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_15_a(Datapath_for_4_ProductSum_for_acc_9_cmp_15_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_15_c(Datapath_for_4_ProductSum_for_acc_9_cmp_15_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_15_z(Datapath_for_4_ProductSum_for_acc_9_cmp_15_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_16_a(Datapath_for_4_ProductSum_for_acc_9_cmp_16_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_16_c(Datapath_for_4_ProductSum_for_acc_9_cmp_16_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_16_z(Datapath_for_4_ProductSum_for_acc_9_cmp_16_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_17_a(Datapath_for_4_ProductSum_for_acc_9_cmp_17_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_17_c(Datapath_for_4_ProductSum_for_acc_9_cmp_17_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_17_z(Datapath_for_4_ProductSum_for_acc_9_cmp_17_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_18_a(Datapath_for_4_ProductSum_for_acc_9_cmp_18_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_18_c(Datapath_for_4_ProductSum_for_acc_9_cmp_18_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_18_z(Datapath_for_4_ProductSum_for_acc_9_cmp_18_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_19_a(Datapath_for_4_ProductSum_for_acc_9_cmp_19_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_19_c(Datapath_for_4_ProductSum_for_acc_9_cmp_19_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_19_z(Datapath_for_4_ProductSum_for_acc_9_cmp_19_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_20_a(Datapath_for_4_ProductSum_for_acc_9_cmp_20_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_20_c(Datapath_for_4_ProductSum_for_acc_9_cmp_20_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_20_z(Datapath_for_4_ProductSum_for_acc_9_cmp_20_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_21_a(Datapath_for_4_ProductSum_for_acc_9_cmp_21_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_21_c(Datapath_for_4_ProductSum_for_acc_9_cmp_21_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_21_z(Datapath_for_4_ProductSum_for_acc_9_cmp_21_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_22_a(Datapath_for_4_ProductSum_for_acc_9_cmp_22_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_22_c(Datapath_for_4_ProductSum_for_acc_9_cmp_22_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_22_z(Datapath_for_4_ProductSum_for_acc_9_cmp_22_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_23_a(Datapath_for_4_ProductSum_for_acc_9_cmp_23_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_23_c(Datapath_for_4_ProductSum_for_acc_9_cmp_23_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_23_z(Datapath_for_4_ProductSum_for_acc_9_cmp_23_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_24_a(Datapath_for_4_ProductSum_for_acc_9_cmp_24_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_24_c(Datapath_for_4_ProductSum_for_acc_9_cmp_24_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_24_z(Datapath_for_4_ProductSum_for_acc_9_cmp_24_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_25_a(Datapath_for_4_ProductSum_for_acc_9_cmp_25_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_25_c(Datapath_for_4_ProductSum_for_acc_9_cmp_25_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_25_z(Datapath_for_4_ProductSum_for_acc_9_cmp_25_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_26_a(Datapath_for_4_ProductSum_for_acc_9_cmp_26_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_26_c(Datapath_for_4_ProductSum_for_acc_9_cmp_26_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_26_z(Datapath_for_4_ProductSum_for_acc_9_cmp_26_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_27_a(Datapath_for_4_ProductSum_for_acc_9_cmp_27_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_27_c(Datapath_for_4_ProductSum_for_acc_9_cmp_27_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_27_z(Datapath_for_4_ProductSum_for_acc_9_cmp_27_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_28_a(Datapath_for_4_ProductSum_for_acc_9_cmp_28_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_28_c(Datapath_for_4_ProductSum_for_acc_9_cmp_28_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_28_z(Datapath_for_4_ProductSum_for_acc_9_cmp_28_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_29_a(Datapath_for_4_ProductSum_for_acc_9_cmp_29_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_29_c(Datapath_for_4_ProductSum_for_acc_9_cmp_29_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_29_z(Datapath_for_4_ProductSum_for_acc_9_cmp_29_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_30_a(Datapath_for_4_ProductSum_for_acc_9_cmp_30_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_30_c(Datapath_for_4_ProductSum_for_acc_9_cmp_30_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_30_z(Datapath_for_4_ProductSum_for_acc_9_cmp_30_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_31_a(Datapath_for_4_ProductSum_for_acc_9_cmp_31_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_31_c(Datapath_for_4_ProductSum_for_acc_9_cmp_31_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_31_z(Datapath_for_4_ProductSum_for_acc_9_cmp_31_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_32_a(Datapath_for_4_ProductSum_for_acc_9_cmp_32_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_32_c(Datapath_for_4_ProductSum_for_acc_9_cmp_32_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_32_z(Datapath_for_4_ProductSum_for_acc_9_cmp_32_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_33_a(Datapath_for_4_ProductSum_for_acc_9_cmp_33_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_33_c(Datapath_for_4_ProductSum_for_acc_9_cmp_33_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_33_z(Datapath_for_4_ProductSum_for_acc_9_cmp_33_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_34_a(Datapath_for_4_ProductSum_for_acc_9_cmp_34_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_34_c(Datapath_for_4_ProductSum_for_acc_9_cmp_34_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_34_z(Datapath_for_4_ProductSum_for_acc_9_cmp_34_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_35_a(Datapath_for_4_ProductSum_for_acc_9_cmp_35_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_35_c(Datapath_for_4_ProductSum_for_acc_9_cmp_35_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_35_z(Datapath_for_4_ProductSum_for_acc_9_cmp_35_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_36_a(Datapath_for_4_ProductSum_for_acc_9_cmp_36_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_36_c(Datapath_for_4_ProductSum_for_acc_9_cmp_36_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_36_z(Datapath_for_4_ProductSum_for_acc_9_cmp_36_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_37_a(Datapath_for_4_ProductSum_for_acc_9_cmp_37_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_37_c(Datapath_for_4_ProductSum_for_acc_9_cmp_37_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_37_z(Datapath_for_4_ProductSum_for_acc_9_cmp_37_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_38_a(Datapath_for_4_ProductSum_for_acc_9_cmp_38_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_38_c(Datapath_for_4_ProductSum_for_acc_9_cmp_38_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_38_z(Datapath_for_4_ProductSum_for_acc_9_cmp_38_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_39_a(Datapath_for_4_ProductSum_for_acc_9_cmp_39_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_39_c(Datapath_for_4_ProductSum_for_acc_9_cmp_39_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_39_z(Datapath_for_4_ProductSum_for_acc_9_cmp_39_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_40_a(Datapath_for_4_ProductSum_for_acc_9_cmp_40_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_40_c(Datapath_for_4_ProductSum_for_acc_9_cmp_40_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_40_z(Datapath_for_4_ProductSum_for_acc_9_cmp_40_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_41_a(Datapath_for_4_ProductSum_for_acc_9_cmp_41_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_41_c(Datapath_for_4_ProductSum_for_acc_9_cmp_41_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_41_z(Datapath_for_4_ProductSum_for_acc_9_cmp_41_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_42_a(Datapath_for_4_ProductSum_for_acc_9_cmp_42_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_42_c(Datapath_for_4_ProductSum_for_acc_9_cmp_42_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_42_z(Datapath_for_4_ProductSum_for_acc_9_cmp_42_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_43_a(Datapath_for_4_ProductSum_for_acc_9_cmp_43_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_43_c(Datapath_for_4_ProductSum_for_acc_9_cmp_43_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_43_z(Datapath_for_4_ProductSum_for_acc_9_cmp_43_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_44_a(Datapath_for_4_ProductSum_for_acc_9_cmp_44_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_44_c(Datapath_for_4_ProductSum_for_acc_9_cmp_44_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_44_z(Datapath_for_4_ProductSum_for_acc_9_cmp_44_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_45_a(Datapath_for_4_ProductSum_for_acc_9_cmp_45_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_45_c(Datapath_for_4_ProductSum_for_acc_9_cmp_45_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_45_z(Datapath_for_4_ProductSum_for_acc_9_cmp_45_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_46_a(Datapath_for_4_ProductSum_for_acc_9_cmp_46_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_46_c(Datapath_for_4_ProductSum_for_acc_9_cmp_46_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_46_z(Datapath_for_4_ProductSum_for_acc_9_cmp_46_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_47_a(Datapath_for_4_ProductSum_for_acc_9_cmp_47_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_47_c(Datapath_for_4_ProductSum_for_acc_9_cmp_47_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_47_z(Datapath_for_4_ProductSum_for_acc_9_cmp_47_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_48_a(Datapath_for_4_ProductSum_for_acc_9_cmp_48_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_48_c(Datapath_for_4_ProductSum_for_acc_9_cmp_48_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_48_z(Datapath_for_4_ProductSum_for_acc_9_cmp_48_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_49_a(Datapath_for_4_ProductSum_for_acc_9_cmp_49_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_49_c(Datapath_for_4_ProductSum_for_acc_9_cmp_49_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_49_z(Datapath_for_4_ProductSum_for_acc_9_cmp_49_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_50_a(Datapath_for_4_ProductSum_for_acc_9_cmp_50_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_50_c(Datapath_for_4_ProductSum_for_acc_9_cmp_50_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_50_z(Datapath_for_4_ProductSum_for_acc_9_cmp_50_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_51_a(Datapath_for_4_ProductSum_for_acc_9_cmp_51_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_51_c(Datapath_for_4_ProductSum_for_acc_9_cmp_51_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_51_z(Datapath_for_4_ProductSum_for_acc_9_cmp_51_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_52_a(Datapath_for_4_ProductSum_for_acc_9_cmp_52_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_52_c(Datapath_for_4_ProductSum_for_acc_9_cmp_52_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_52_z(Datapath_for_4_ProductSum_for_acc_9_cmp_52_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_53_a(Datapath_for_4_ProductSum_for_acc_9_cmp_53_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_53_c(Datapath_for_4_ProductSum_for_acc_9_cmp_53_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_53_z(Datapath_for_4_ProductSum_for_acc_9_cmp_53_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_54_a(Datapath_for_4_ProductSum_for_acc_9_cmp_54_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_54_c(Datapath_for_4_ProductSum_for_acc_9_cmp_54_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_54_z(Datapath_for_4_ProductSum_for_acc_9_cmp_54_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_55_a(Datapath_for_4_ProductSum_for_acc_9_cmp_55_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_55_c(Datapath_for_4_ProductSum_for_acc_9_cmp_55_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_55_z(Datapath_for_4_ProductSum_for_acc_9_cmp_55_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_56_a(Datapath_for_4_ProductSum_for_acc_9_cmp_56_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_56_c(Datapath_for_4_ProductSum_for_acc_9_cmp_56_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_56_z(Datapath_for_4_ProductSum_for_acc_9_cmp_56_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_57_a(Datapath_for_4_ProductSum_for_acc_9_cmp_57_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_57_c(Datapath_for_4_ProductSum_for_acc_9_cmp_57_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_57_z(Datapath_for_4_ProductSum_for_acc_9_cmp_57_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_58_a(Datapath_for_4_ProductSum_for_acc_9_cmp_58_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_58_c(Datapath_for_4_ProductSum_for_acc_9_cmp_58_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_58_z(Datapath_for_4_ProductSum_for_acc_9_cmp_58_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_59_a(Datapath_for_4_ProductSum_for_acc_9_cmp_59_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_59_c(Datapath_for_4_ProductSum_for_acc_9_cmp_59_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_59_z(Datapath_for_4_ProductSum_for_acc_9_cmp_59_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_60_a(Datapath_for_4_ProductSum_for_acc_9_cmp_60_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_60_c(Datapath_for_4_ProductSum_for_acc_9_cmp_60_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_60_z(Datapath_for_4_ProductSum_for_acc_9_cmp_60_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_61_a(Datapath_for_4_ProductSum_for_acc_9_cmp_61_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_61_c(Datapath_for_4_ProductSum_for_acc_9_cmp_61_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_61_z(Datapath_for_4_ProductSum_for_acc_9_cmp_61_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_62_a(Datapath_for_4_ProductSum_for_acc_9_cmp_62_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_62_c(Datapath_for_4_ProductSum_for_acc_9_cmp_62_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_62_z(Datapath_for_4_ProductSum_for_acc_9_cmp_62_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_63_a(Datapath_for_4_ProductSum_for_acc_9_cmp_63_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_63_c(Datapath_for_4_ProductSum_for_acc_9_cmp_63_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_63_z(Datapath_for_4_ProductSum_for_acc_9_cmp_63_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_1_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_1_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_2_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_2_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_3_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_3_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_4_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_4_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_5_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_5_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_6_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_6_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_7_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_7_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_41_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_41_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_41_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_41_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_42_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_42_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_42_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_42_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_43_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_43_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_43_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_43_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_44_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_44_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_44_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_44_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_45_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_45_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_45_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_45_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_46_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_46_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_46_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_46_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_47_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_47_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_47_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_47_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff)
    );
endmodule



