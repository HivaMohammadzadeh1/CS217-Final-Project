
//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 02:51:36 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [168:0] this_dat;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [127:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_dat[127:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_dat[151:128];
  wire  nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_dat[168];
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd128)) data_data_rsci (
      .d(nl_data_data_rsci_d[127:0]),
      .z(data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d),
      .z(data_rw_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd154),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [168:0] this_dat;
  output [127:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 04:38:56 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [137:0] this_dat;
  output [127:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [127:0] nl_data_data_data_rsci_d;
  assign nl_data_data_data_rsci_d = this_dat[127:0];
  wire [7:0] nl_data_logical_addr_rsci_d;
  assign nl_data_logical_addr_rsci_d = this_dat[137:130];
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd7),
  .width(32'sd128)) data_data_data_rsci (
      .d(nl_data_data_data_rsci_d[127:0]),
      .z(data_data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd9),
  .width(32'sd8)) data_logical_addr_rsci (
      .d(nl_data_logical_addr_rsci_d[7:0]),
      .z(data_logical_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd11),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd153),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [137:0] this_dat;
  output [127:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_data_rsc_z(data_data_data_rsc_z),
      .data_logical_addr_rsc_z(data_logical_addr_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 04:38:53 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [255:0] this_dat;
  reg [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [255:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd13),
  .width(32'sd256)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd152),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd156)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 01:32:50 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd15),
  .width(32'sd1)) data_rsci (
      .d(this_dat),
      .z(data_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd17),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd151),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 02:51:33 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [127:0] this_dat;
  reg [127:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [127:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd18),
  .width(32'sd128)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd150),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd155)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [127:0] this_dat;
  input [127:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module PECore_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // spyglass disable SYNTH_5121,W240
    input                s_rst;  // spyglass disable SYNTH_5121,W240
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a; //spyglass disable FlopEConst
                b_reg[0] <= b; //spyglass disable FlopEConst
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> ./PECore_mgc_muladd1_beh.v 
//muladd1
module PECore_mgc_muladd1(a,b,c,cst,d,z);
  // operation is z = a * (b + d) + c + cst
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_cst = 0;
  parameter signd_cst = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_axb = 1;
  parameter add_c = 1;
  parameter add_d = 1;
  parameter use_const = 1;

  function integer is_square_op;
    input integer alen;
  begin
    if (alen > 1) is_square_op = 0;
    else       is_square_op = 1;
  end endfunction

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_cst-1:0] cst; // spyglass disable SYNTH_5121,W240
  input  [width_d-1:0] d;
  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa;
  reg [width_b-signd_b:0] bb;
  reg [width_c-signd_c:0] cc;
  reg [width_d-signd_d:0] dd;
  reg [width_cst-signd_cst:0] cstin;

  localparam width_bd = (width_d) ? 1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b
                                                                          : width_d - signd_d)
                                  : width_b - signd_b;
  localparam is_square = is_square_op(width_a);
  localparam axb_len = (is_square)?width_bd+1+width_bd+1:width_a-signd_a+1+width_bd+1;

  reg [width_bd:0] bd;
  reg [axb_len-1:0] axb;



  // make all inputs signed
  always @(*) aa = signd_a ? a : {1'b0, a};
  always @(*) bb = signd_b ? b : {1'b0, b};
  generate if (width_c != 0) begin
    always @(*) cc = signd_c ? c : {1'b0, c};
  end endgenerate

  generate if (width_d) begin
    if ( !is_square) begin
      (* keep ="true" *) reg [width_d-signd_d:0] d_keep;
      always @(*) d_keep = signd_d ? d : {1'b0, d};
      always @(*) dd = d_keep;
    end else begin
      always @(*) dd = signd_d ? d : {1'b0, d};
    end
  end endgenerate

  always @(*) cstin = signd_cst ? cst : {1'b0, cst};

  // perform pre-adder
  generate
    if (width_d != 0) begin
      if (add_d) begin always @(*)  bd = $signed(bb) + $signed(dd); end
      else       begin always @(*)  bd = $signed(bb) - $signed(dd); end
    end else     begin always @(*)  bd = $signed(bb); end
  endgenerate

  generate
    if (is_square)
      always @(*) axb = $signed(bd) * $signed(bd);
    else
      always @(*) axb = $signed(aa) * $signed(bd);
  endgenerate

  // perform muladd1
  wire [width_z-1:0]  zz;

  generate
    if (use_const) begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc) + $signed(cstin); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc) + $signed(cstin); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb) + $signed(cstin); end else
      if (!add_axb && !add_c && width_c) begin assign zz = $signed(cstin) - $signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb) + $signed(cstin); end else
                                         begin assign zz = $signed(cstin) - $signed(axb); end
    end  else begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb); end else
      if (!add_axb && !add_c && width_c) begin assign zz = -$signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb); end else
                                         begin assign zz = -$signed(axb); end
    end
  endgenerate

  // adjust output
  assign z = zz;
endmodule // mgc_muladd1

//------> ./PECore_mgc_shift_l_beh_v5.v 
module PECore_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./PECore_mgc_mul2add1_pipe_beh.v 
//muladd1
module PECore_mgc_mul2add1_pipe(a,b,b2,c,d,d2,cst,clk,en,a_rst,s_rst,z);
  parameter gentype = 0;
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_b2 = 0;
  parameter signd_b2 = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_d2 = 0;
  parameter signd_d2 = 0;
  parameter width_e = 0;
  parameter signd_e = 0;
  parameter width_z = 0;
  parameter isadd = 1;
  parameter add_b2 = 1;
  parameter add_d2 = 1;
  parameter use_const = 1;
  parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
  parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
  parameter    a_rst_active =  1'b1;  // unused
  parameter    s_rst_active =  1'b1;  // unused
  parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
  parameter integer n_inreg = 32'd0;  // number of input registers

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_b2-1:0] b2; // spyglass disable SYNTH_5121,W240
  input  [width_c-1:0] c;
  input  [width_d-1:0] d;
  input  [width_d2-1:0] d2; // spyglass disable SYNTH_5121,W240
  input  [width_e-1:0] cst; // spyglass disable SYNTH_5121,W240

  input                clk;    // clock
  input                en;     // enable
  input                a_rst;  // spyglass disable SYNTH_5121,W240
  input                s_rst;  // spyglass disable SYNTH_5121,W240

  output [width_z-1:0] z;

  function integer MIN;
    input integer a, b;
  begin
    if (a > b) MIN = b;
    else       MIN = a;
  end endfunction

  function integer f_axb_stages;
    input integer gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d;
  begin
    if (gentype%2==0) begin
      if ((n_inreg > 1) && (width_a>18 | width_b>=19+signd_b | width_c>18 | width_d>=19+signd_d ))
        f_axb_stages = 1;
      else
        f_axb_stages = 0;
    end else begin
      if (n_inreg>1)
        f_axb_stages = 1;
      else
        f_axb_stages = 0;
    end
  end endfunction

  function integer f_cxd_stages;
    input integer gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d;
  begin
    if (gentype%2==0) begin
      f_cxd_stages = 0;
    end else begin
      if (n_inreg>1)
        f_cxd_stages = MIN(n_inreg-1,3);
      else
        f_cxd_stages = 0;
    end
  end endfunction

  function integer f_preadd_stages;
    input integer gentype,n_inreg,width_preaddin;
  begin
    if (gentype%2==0) begin
      f_preadd_stages = 0;
    end else begin
      if (n_inreg>1) begin
        if (width_preaddin>0)
          f_preadd_stages = 1;
        else
          f_preadd_stages = 0;
      end else
        f_preadd_stages = 0;
    end
  end endfunction

  function integer MAX;
    input integer LEFT, RIGHT;
  begin
    if (LEFT > RIGHT) MAX = LEFT;
    else              MAX = RIGHT;
  end endfunction

  function integer PREADDLEN;
    input integer b_len, d_len, width_d;
  begin
    if(width_d>0) PREADDLEN = MAX(b_len,d_len) + 1;
    else        PREADDLEN = b_len;
  end endfunction
  function integer PREADDMULLEN;
    input integer a_len, b_len, d_len, width_d;
  begin
    PREADDMULLEN = a_len + PREADDLEN(b_len,d_len,width_d);
  end endfunction

  localparam axb_stages = f_axb_stages(gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d);
  localparam cxd_stages = f_cxd_stages(gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d);
  localparam preadd_ab_stages = f_preadd_stages(gentype, n_inreg - axb_stages,width_b2);
  localparam preadd_cd_stages = f_preadd_stages(gentype, n_inreg - cxd_stages,width_d2);
  localparam e_stages  = (use_const>1)?n_inreg:0;
  localparam a_stages  = n_inreg - axb_stages;
  localparam b_stages  = n_inreg - axb_stages - preadd_ab_stages;
  localparam c_stages  = n_inreg - cxd_stages;
  localparam d_stages  = n_inreg - cxd_stages - preadd_cd_stages;
  localparam b2_stages  = (width_b2>0)?b_stages:0;
  localparam d2_stages  = (width_d2>0)?d_stages:0;

  localparam a_len    = width_a-signd_a+1;
  localparam b_len    = width_b-signd_b+1;
  localparam b2_len   = width_b2-signd_b2+1;
  localparam c_len    = width_c-signd_c+1;
  localparam d_len    = width_d-signd_d+1;
  localparam d2_len   = width_d2-signd_d2+1;
  localparam e_len    = width_e-signd_e+1;
  localparam bb2_len  = PREADDLEN(b_len, b2_len, width_b2);
  localparam dd2_len  = PREADDLEN(d_len, d2_len, width_d2);
  localparam axb_len  = PREADDMULLEN(a_len, b_len, b2_len, width_b2);
  localparam cxd_len  = PREADDMULLEN(c_len, d_len, d2_len, width_d2);
  localparam z_len    = width_z;

  reg [a_len-1:0]  aa  [a_stages:0];
  reg [b_len-1:0]  bb  [b_stages:0];
  reg [b2_len-1:0] bb2 [b2_stages:0];
  reg [c_len-1:0]  cc  [c_stages:0];
  reg [d_len-1:0]  dd  [d_stages:0];
  reg [d2_len-1:0] dd2 [d2_stages:0];
  reg [e_len-1:0]  ee  [e_stages:0];



  genvar i;

  // make all inputs signed
  always @(*) aa[a_stages] = signd_a ? a : {1'b0, a}; //spyglass disable W164a W164b
  always @(*) bb[b_stages] = signd_b ? b : {1'b0, b}; //spyglass disable W164a W164b
  generate if (width_b2>0) begin
    (* keep ="true" *) reg [b2_len-1:0] b2_keep;
    always @(*) b2_keep = signd_b2 ? b2 : {1'b0, b2}; //spyglass disable W164a W164b
    always @(*) bb2[b2_stages] = b2_keep;
  end endgenerate
  always @(*) cc[c_stages] = signd_c ? c : {1'b0, c}; //spyglass disable W164a W164b
  always @(*) dd[d_stages] = signd_d ? d : {1'b0, d}; //spyglass disable W164a W164b
  generate if (width_d2>0) begin
    (* keep ="true" *) reg [d2_len-1:0] d2_keep;
    always @(*) d2_keep = signd_d2 ? d2 : {1'b0, d2}; //spyglass disable W164a W164b
    always @(*) dd2[d2_stages] = d2_keep;
  end endgenerate

  generate if (use_const>0) begin
    always @(*) ee[e_stages] = signd_e ? cst : {1'b0, cst}; //spyglass disable W164a W164b

    // input registers
    if (e_stages>0) begin
    for(i = e_stages-1; i >= 0; i=i-1) begin:in_pipe_e
      if (clock_edge == 1'b1) begin:pos
        always @(posedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
      end else begin:neg
        always @(negedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
      end
    end end
  end endgenerate
  generate if (a_stages>0) begin
  for(i = a_stages-1; i >= 0; i=i-1) begin:in_pipe_a
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (b_stages>0) begin
  for(i = b_stages-1; i >= 0; i=i-1) begin:in_pipe_b
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];
    end
  end end endgenerate
  generate if (c_stages>0) begin
  for(i = c_stages-1; i >= 0; i=i-1) begin:in_pipe_c
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (d_stages>0) begin
  for(i = d_stages-1; i >= 0; i=i-1) begin:in_pipe_d
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) dd[i] <= dd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) dd[i] <= dd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (b2_stages>0) begin
  for(i = b2_stages-1; i >= 0; i=i-1) begin:in_pipe_b2
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb2[i] <= bb2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb2[i] <= bb2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (d2_stages>0) begin
  for(i = d2_stages-1; i >= 0; i=i-1) begin:in_pipe_d2
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) dd2[i] <= dd2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) dd2[i] <= dd2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg [bb2_len-1:0] b_bb2[preadd_ab_stages:0];
  reg [dd2_len-1:0] d_dd2[preadd_cd_stages:0];

  //perform first preadd
  generate
    if (width_b2>0) begin
      if (add_b2) begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]) + $signed(bb2[0]); end
      else        begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]) - $signed(bb2[0]); end
    end else      begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]); end
  endgenerate
  generate if (preadd_ab_stages>0) begin
  for(i = preadd_ab_stages-1; i >= 0; i=i-1) begin:preaddab_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) b_bb2[i] <= b_bb2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) b_bb2[i] <= b_bb2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  //perform second preadd
  generate
    if (width_d2>0) begin
      if (add_d2) begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]) + $signed(dd2[0]); end
      else        begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]) - $signed(dd2[0]); end
    end else      begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]); end
  endgenerate
  generate if (preadd_cd_stages>0) begin
  for(i = preadd_cd_stages-1; i >= 0; i=i-1) begin:preaddcd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) d_dd2[i] <= d_dd2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) d_dd2[i] <= d_dd2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // perform first multiplication
  reg [axb_len-1:0] axb[axb_stages:0];

  always @(*) axb[axb_stages] = $signed(aa[0]) * $signed(b_bb2[0]);
  generate if (axb_stages>0) begin
  for(i = axb_stages-1; i >= 0; i=i-1) begin:axb_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];
    end
  end end endgenerate

  // perform second multiplication
  reg [cxd_len-1:0] cxd[cxd_stages:0];

  always @(*) cxd[cxd_stages] = $signed(cc[0]) * $signed(d_dd2[0]);
  generate if (cxd_stages>0) begin
  for(i = cxd_stages-1; i >= 0; i=i-1) begin:cxd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cxd[i] <= cxd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cxd[i] <= cxd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg [z_len-1:0]  zz[stages-1:0];
  generate
    if (use_const>1) begin
      reg [z_len-1:0] aux_val;
      if ( isadd) begin
        always @(*) aux_val = $signed(axb[0]) + $signed(cxd[0]);
      end else begin
        always @(*) aux_val = $signed(axb[0]) - $signed(cxd[0]);
      end
      always @(*) zz[stages-1] = $signed(ee[0]) + $signed(aux_val) ;
    end else begin
      if (use_const>0) begin
        if ( isadd) begin always @(*) zz[stages-1] = $signed(axb[0]) + $signed(cxd[0]) + $signed(ee[0]); end else
                    begin always @(*) zz[stages-1] = $signed(axb[0]) - $signed(cxd[0]) + $signed(ee[0]); end
      end else begin
        if ( isadd) begin always @(*) zz[stages-1] = $signed(axb[0]) + $signed(cxd[0]); end else
                    begin always @(*) zz[stages-1] = $signed(axb[0]) - $signed(cxd[0]); end
      end
    end
  endgenerate

  // Output registers:
  generate if (stages>1) begin
  for(i = stages-2; i >= 0; i=i-1) begin:out_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // adjust output
  assign z = zz[0];
endmodule // mgc_mul2add1_pipe

//------> /cad/mentor/2024.2_1/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)
// suppress_sim_read_addr_range_errs:  0 - report errors  1 - suppress errors

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 ,
  parameter suppress_sim_read_addr_range_errs = 1 
  
)( clk,clken,d,q,radr,re,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input  re;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" , syn_ramstyle = "block" *)
  reg [data_width-1:0] mem [depth-1:0];
  integer j;
  initial for (j = 0; j < depth; j = j + 1) mem[j] = 0;
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr READ_ENABLE re
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg re_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
          re_reg <= re;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./PECore.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 04:51:42 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_128_4096_1_4096_128_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_128_4096_1_4096_128_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [127:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [127:0] d;
  output [11:0] wadr;
  input clken_d;
  input [127:0] d_d;
  output [127:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_PECoreRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_PECoreRun_fsm (
  clk, rst, PECoreRun_wen, fsm_output
);
  input clk;
  input rst;
  input PECoreRun_wen;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for PECore_PECore_PECoreRun_PECoreRun_fsm_1
  parameter
    PECoreRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : PECore_PECore_PECoreRun_PECoreRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // PECoreRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= PECoreRun_rlp_C_0;
    end
    else if ( PECoreRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_staller
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_staller (
  clk, rst, PECoreRun_wen, PECoreRun_wten, act_port_Push_mioi_wen_comp, rva_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PECoreRun_wen;
  output PECoreRun_wten;
  input act_port_Push_mioi_wen_comp;
  input rva_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg PECoreRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign PECoreRun_wen = act_port_Push_mioi_wen_comp & rva_out_Push_mioi_wen_comp;
  assign PECoreRun_wten = PECoreRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECoreRun_wten_reg <= 1'b0;
    end
    else begin
      PECoreRun_wten_reg <= ~ PECoreRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_wait_dp (
  weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      Datapath_for_4_ProductSum_for_acc_5_cmp_en, Datapath_for_4_ProductSum_for_acc_5_cmp_5_en,
      PECoreRun_wen, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg,
      PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo, PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg,
      PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en, PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_1,
      PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg_1, PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en,
      Datapath_for_4_ProductSum_for_acc_5_cmp_cgo, Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg,
      Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_5, Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg_5
);
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output Datapath_for_4_ProductSum_for_acc_5_cmp_en;
  output Datapath_for_4_ProductSum_for_acc_5_cmp_5_en;
  input PECoreRun_wen;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg;
  input PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo;
  input PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg;
  output PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en;
  input PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_1;
  input PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg_1;
  output PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en;
  input Datapath_for_4_ProductSum_for_acc_5_cmp_cgo;
  input Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg;
  input Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_5;
  input Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg_5;



  // Interconnect Declarations for Component Instantiations 
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg);
  assign PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en = PECoreRun_wen & (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo
      | PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg);
  assign PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en = PECoreRun_wen & (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_1
      | PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg_1);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_en = ~(PECoreRun_wen & (Datapath_for_4_ProductSum_for_acc_5_cmp_cgo
      | Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg));
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_5_en = ~(PECoreRun_wen & (Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_5
      | Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg_5));
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  PECoreRun_wen, rva_out_Push_mioi_oswt, rva_out_Push_mioi_biwt, rva_out_Push_mioi_bdwt,
      rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & PECoreRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt)
      & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & rva_out_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt,
      start_PopNB_mioi_biwt_pff, start_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_biwt_pff;
  input start_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & PECoreRun_wen;
  assign start_PopNB_mioi_biwt = (~ PECoreRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_biwt_pff = PECoreRun_wen & start_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp (
  clk, rst, act_port_Push_mioi_oswt, act_port_Push_mioi_wen_comp, act_port_Push_mioi_biwt,
      act_port_Push_mioi_bdwt, act_port_Push_mioi_bcwt
);
  input clk;
  input rst;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input act_port_Push_mioi_biwt;
  input act_port_Push_mioi_bdwt;
  output act_port_Push_mioi_bcwt;
  reg act_port_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_wen_comp = (~ act_port_Push_mioi_oswt) | act_port_Push_mioi_biwt
      | act_port_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_Push_mioi_bcwt <= ~((~(act_port_Push_mioi_bcwt | act_port_Push_mioi_biwt))
          | act_port_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl (
  PECoreRun_wen, act_port_Push_mioi_oswt, act_port_Push_mioi_biwt, act_port_Push_mioi_bdwt,
      act_port_Push_mioi_bcwt, act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      act_port_Push_mioi_ccs_ccore_done_sync_vld, act_port_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_biwt;
  output act_port_Push_mioi_bdwt;
  input act_port_Push_mioi_bcwt;
  output act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input act_port_Push_mioi_ccs_ccore_done_sync_vld;
  input act_port_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_bdwt = act_port_Push_mioi_oswt & PECoreRun_wen;
  assign act_port_Push_mioi_biwt = act_port_Push_mioi_oswt & (~ act_port_Push_mioi_bcwt)
      & act_port_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & act_port_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
    (
  clk, rst, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt,
      input_port_PopNB_mioi_return_rsc_z_mxwt, input_port_PopNB_mioi_biwt, input_port_PopNB_mioi_bdwt,
      input_port_PopNB_mioi_data_data_data_rsc_z, input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_biwt;
  input input_port_PopNB_mioi_bdwt;
  input [127:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  input [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  input input_port_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg input_port_PopNB_mioi_bcwt;
  reg [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_bfwt;
  reg [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt;
  reg input_port_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_data_data_data_rsc_z_mxwt = MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z,
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt = MUX_v_8_2_2(input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z,
      input_port_PopNB_mioi_return_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      input_port_PopNB_mioi_bcwt <= ~((~(input_port_PopNB_mioi_bcwt | input_port_PopNB_mioi_biwt))
          | input_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= 8'b00000000;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( input_port_PopNB_mioi_biwt ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= input_port_PopNB_mioi_data_data_data_rsc_z;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= input_port_PopNB_mioi_data_logical_addr_rsc_z;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= input_port_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
    (
  PECoreRun_wen, PECoreRun_wten, input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_biwt,
      input_port_PopNB_mioi_bdwt, input_port_PopNB_mioi_biwt_pff, input_port_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output input_port_PopNB_mioi_biwt;
  output input_port_PopNB_mioi_bdwt;
  output input_port_PopNB_mioi_biwt_pff;
  input input_port_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_bdwt = input_port_PopNB_mioi_oswt & PECoreRun_wen;
  assign input_port_PopNB_mioi_biwt = (~ PECoreRun_wten) & input_port_PopNB_mioi_oswt;
  assign input_port_PopNB_mioi_biwt_pff = PECoreRun_wen & input_port_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [127:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  reg [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_128_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_20_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4, rva_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= 20'b00000000000000000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & PECoreRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ PECoreRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = PECoreRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, PECoreRun_wen, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_PECoreRun, rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [127:0] rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_oswt_pff(rva_out_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi (
  clk, rst, start_vld, start_rdy, start_dat, PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_vld(start_vld),
      .this_rdy(start_rdy),
      .this_dat(start_dat),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_biwt_pff(start_PopNB_mioi_biwt_iff),
      .start_PopNB_mioi_oswt_pff(start_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi (
  clk, rst, act_port_vld, act_port_rdy, act_port_dat, PECoreRun_wen, act_port_Push_mioi_oswt,
      act_port_Push_mioi_wen_comp, act_port_Push_mioi_m_data_rsc_dat_PECoreRun, act_port_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input [255:0] act_port_Push_mioi_m_data_rsc_dat_PECoreRun;
  input act_port_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_port_Push_mioi_biwt;
  wire act_port_Push_mioi_bdwt;
  wire act_port_Push_mioi_bcwt;
  wire act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire act_port_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push  act_port_Push_mioi
      (
      .this_vld(act_port_vld),
      .this_rdy(act_port_rdy),
      .this_dat(act_port_dat),
      .m_data_rsc_dat(act_port_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt),
      .act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .act_port_Push_mioi_ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .act_port_Push_mioi_oswt_pff(act_port_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi (
  clk, rst, input_port_vld, input_port_rdy, input_port_dat, PECoreRun_wen, PECoreRun_wten,
      input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt, input_port_PopNB_mioi_return_rsc_z_mxwt,
      input_port_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input input_port_vld;
  output input_port_rdy;
  input [137:0] input_port_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_port_PopNB_mioi_biwt;
  wire input_port_PopNB_mioi_bdwt;
  wire [127:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  wire input_port_PopNB_mioi_return_rsc_z;
  wire input_port_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB  input_port_PopNB_mioi
      (
      .this_vld(input_port_vld),
      .this_rdy(input_port_rdy),
      .this_dat(input_port_dat),
      .data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .return_rsc_z(input_port_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(input_port_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(input_port_PopNB_mioi_oswt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_biwt_pff(input_port_PopNB_mioi_biwt_iff),
      .input_port_PopNB_mioi_oswt_pff(input_port_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .input_port_PopNB_mioi_return_rsc_z(input_port_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt,
      rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG, weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d, Datapath_for_4_ProductSum_for_acc_5_cmp_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_c, Datapath_for_4_ProductSum_for_acc_5_cmp_en,
      Datapath_for_4_ProductSum_for_acc_5_cmp_z, Datapath_for_4_ProductSum_for_acc_5_cmp_1_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_1_c, Datapath_for_4_ProductSum_for_acc_5_cmp_1_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_2_a, Datapath_for_4_ProductSum_for_acc_5_cmp_2_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_2_z, Datapath_for_4_ProductSum_for_acc_5_cmp_3_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_3_c, Datapath_for_4_ProductSum_for_acc_5_cmp_3_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_4_a, Datapath_for_4_ProductSum_for_acc_5_cmp_4_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_4_z, Datapath_for_4_ProductSum_for_acc_5_cmp_5_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_5_c, Datapath_for_4_ProductSum_for_acc_5_cmp_5_en,
      Datapath_for_4_ProductSum_for_acc_5_cmp_5_z, Datapath_for_4_ProductSum_for_acc_5_cmp_6_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_c, Datapath_for_4_ProductSum_for_acc_5_cmp_6_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_7_a, Datapath_for_4_ProductSum_for_acc_5_cmp_7_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_7_z, Datapath_for_4_ProductSum_for_acc_5_cmp_8_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_8_c, Datapath_for_4_ProductSum_for_acc_5_cmp_8_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_9_a, Datapath_for_4_ProductSum_for_acc_5_cmp_9_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_9_z, Datapath_for_4_ProductSum_for_acc_5_cmp_10_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_10_c, Datapath_for_4_ProductSum_for_acc_5_cmp_10_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_11_a, Datapath_for_4_ProductSum_for_acc_5_cmp_11_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_11_z, Datapath_for_4_ProductSum_for_acc_5_cmp_12_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_12_c, Datapath_for_4_ProductSum_for_acc_5_cmp_12_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_13_a, Datapath_for_4_ProductSum_for_acc_5_cmp_13_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_13_z, Datapath_for_4_ProductSum_for_acc_5_cmp_14_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_14_c, Datapath_for_4_ProductSum_for_acc_5_cmp_14_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_15_a, Datapath_for_4_ProductSum_for_acc_5_cmp_15_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_15_z, Datapath_for_4_ProductSum_for_acc_5_cmp_16_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_16_c, Datapath_for_4_ProductSum_for_acc_5_cmp_16_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_17_a, Datapath_for_4_ProductSum_for_acc_5_cmp_17_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_17_z, Datapath_for_4_ProductSum_for_acc_5_cmp_18_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_18_c, Datapath_for_4_ProductSum_for_acc_5_cmp_18_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_19_a, Datapath_for_4_ProductSum_for_acc_5_cmp_19_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_19_z, Datapath_for_4_ProductSum_for_acc_5_cmp_20_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_20_c, Datapath_for_4_ProductSum_for_acc_5_cmp_20_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_21_a, Datapath_for_4_ProductSum_for_acc_5_cmp_21_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_21_z, Datapath_for_4_ProductSum_for_acc_5_cmp_22_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_22_c, Datapath_for_4_ProductSum_for_acc_5_cmp_22_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_23_a, Datapath_for_4_ProductSum_for_acc_5_cmp_23_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_23_z, Datapath_for_4_ProductSum_for_acc_5_cmp_24_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_24_c, Datapath_for_4_ProductSum_for_acc_5_cmp_24_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_25_a, Datapath_for_4_ProductSum_for_acc_5_cmp_25_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_25_z, Datapath_for_4_ProductSum_for_acc_5_cmp_26_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_26_c, Datapath_for_4_ProductSum_for_acc_5_cmp_26_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_27_a, Datapath_for_4_ProductSum_for_acc_5_cmp_27_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_27_z, Datapath_for_4_ProductSum_for_acc_5_cmp_28_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_28_c, Datapath_for_4_ProductSum_for_acc_5_cmp_28_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_29_a, Datapath_for_4_ProductSum_for_acc_5_cmp_29_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_29_z, Datapath_for_4_ProductSum_for_acc_5_cmp_30_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_30_c, Datapath_for_4_ProductSum_for_acc_5_cmp_30_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_31_a, Datapath_for_4_ProductSum_for_acc_5_cmp_31_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_31_z, Datapath_for_4_ProductSum_for_acc_5_cmp_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff, weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [137:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  input [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_c;
  output Datapath_for_4_ProductSum_for_acc_5_cmp_en;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_c;
  output Datapath_for_4_ProductSum_for_acc_5_cmp_5_en;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff;


  // Interconnect Declarations
  wire PECoreRun_wen;
  wire PECoreRun_wten;
  wire [127:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [127:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  wire input_port_PopNB_mioi_return_rsc_z_mxwt;
  wire act_port_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_z;
  wire PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_z;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
  wire fsm_output;
  wire pe_config_UpdateManagerCounter_if_if_unequal_tmp;
  wire [7:0] weight_mem_write_arbxbar_xbar_for_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_7_false_1_operator_7_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_7_false_1_operator_7_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  wire nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_1_tmp;
  wire nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp;
  wire while_mux_1331_tmp;
  wire while_mux_1330_tmp;
  wire while_mux_1329_tmp;
  wire while_mux_1328_tmp;
  wire while_mux_1327_tmp;
  wire while_mux_1326_tmp;
  wire while_mux_1325_tmp;
  wire while_mux_1324_tmp;
  wire while_mux_1323_tmp;
  wire while_mux_1322_tmp;
  wire while_mux_1321_tmp;
  wire while_mux_1320_tmp;
  wire while_mux_1319_tmp;
  wire while_mux_1318_tmp;
  wire while_mux_1283_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_125_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_5_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_8_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp;
  wire weight_mem_run_3_for_weight_mem_run_3_for_and_3_tmp;
  wire while_and_30_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  wire and_dcpl_6;
  wire and_dcpl_7;
  wire and_dcpl_10;
  wire and_dcpl_28;
  wire and_dcpl_35;
  wire and_dcpl_41;
  wire and_dcpl_45;
  wire and_dcpl_48;
  wire mux_tmp;
  wire and_dcpl_59;
  wire and_dcpl_71;
  wire and_dcpl_78;
  wire and_dcpl_80;
  wire and_dcpl_82;
  wire or_dcpl_28;
  wire or_dcpl_31;
  wire and_dcpl_84;
  wire and_dcpl_86;
  wire or_dcpl_35;
  wire and_dcpl_88;
  wire or_dcpl_42;
  wire and_dcpl_90;
  wire or_dcpl_52;
  wire and_dcpl_92;
  wire or_dcpl_53;
  wire or_dcpl_59;
  wire and_dcpl_94;
  wire or_dcpl_60;
  wire or_dcpl_63;
  wire or_dcpl_64;
  wire and_dcpl_136;
  wire and_dcpl_137;
  wire and_dcpl_138;
  wire and_dcpl_139;
  wire and_dcpl_140;
  wire and_dcpl_141;
  wire and_dcpl_142;
  wire and_dcpl_143;
  wire and_dcpl_144;
  wire and_dcpl_146;
  wire and_dcpl_154;
  wire mux_tmp_13;
  wire or_tmp_27;
  wire or_tmp_28;
  wire mux_tmp_14;
  wire mux_tmp_15;
  wire mux_tmp_16;
  wire mux_tmp_18;
  wire mux_tmp_27;
  wire and_dcpl_167;
  wire and_dcpl_168;
  wire and_dcpl_169;
  wire and_dcpl_170;
  wire and_dcpl_172;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_179;
  wire and_dcpl_180;
  wire and_dcpl_182;
  wire and_dcpl_183;
  wire and_dcpl_185;
  wire and_dcpl_186;
  wire and_dcpl_189;
  wire and_dcpl_193;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire or_dcpl_132;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire and_dcpl_207;
  wire and_dcpl_208;
  wire and_dcpl_210;
  wire and_dcpl_212;
  wire and_dcpl_216;
  wire and_dcpl_220;
  wire mux_tmp_41;
  wire mux_tmp_42;
  wire mux_tmp_44;
  wire and_dcpl_237;
  wire and_dcpl_238;
  wire and_dcpl_241;
  wire and_dcpl_252;
  wire or_tmp_54;
  wire not_tmp_147;
  wire mux_tmp_56;
  wire and_dcpl_265;
  wire and_dcpl_266;
  wire or_tmp_59;
  wire or_tmp_60;
  wire mux_tmp_65;
  wire or_tmp_61;
  wire mux_tmp_67;
  wire or_tmp_63;
  wire mux_tmp_75;
  wire or_tmp_67;
  wire mux_tmp_76;
  wire and_dcpl_279;
  wire and_dcpl_292;
  wire and_dcpl_297;
  wire and_dcpl_325;
  wire and_dcpl_354;
  wire and_dcpl_362;
  wire and_dcpl_365;
  wire and_dcpl_379;
  wire and_dcpl_393;
  wire and_dcpl_400;
  wire and_dcpl_438;
  wire and_dcpl_443;
  wire or_dcpl_198;
  wire and_dcpl_461;
  wire and_dcpl_468;
  wire and_dcpl_481;
  wire and_dcpl_482;
  wire mux_tmp_92;
  wire and_dcpl_488;
  wire and_dcpl_523;
  wire and_dcpl_527;
  wire or_tmp_79;
  wire and_dcpl_536;
  wire nor_tmp_17;
  wire not_tmp_249;
  wire and_dcpl_538;
  wire not_tmp_252;
  wire mux_tmp_102;
  wire and_tmp;
  wire and_tmp_1;
  wire or_tmp_105;
  wire and_tmp_2;
  wire or_tmp_109;
  wire and_tmp_3;
  wire and_tmp_4;
  wire mux_tmp_118;
  wire and_tmp_5;
  wire or_tmp_121;
  wire nand_tmp_1;
  wire or_tmp_123;
  wire or_tmp_129;
  wire and_dcpl_561;
  wire or_dcpl_219;
  wire or_dcpl_222;
  wire and_dcpl_579;
  wire and_dcpl_580;
  wire and_dcpl_582;
  wire or_dcpl_225;
  wire and_dcpl_614;
  wire and_dcpl_618;
  wire or_dcpl_226;
  wire or_dcpl_231;
  wire or_dcpl_233;
  wire and_dcpl_625;
  wire and_dcpl_636;
  wire or_dcpl_273;
  wire and_dcpl_639;
  wire and_dcpl_643;
  wire or_dcpl_277;
  wire and_dcpl_652;
  wire and_dcpl_655;
  wire and_dcpl_665;
  wire and_dcpl_666;
  wire or_dcpl_279;
  wire nor_tmp_38;
  wire or_tmp_138;
  wire or_tmp_139;
  wire nor_tmp_41;
  wire or_tmp_140;
  wire or_tmp_141;
  wire mux_tmp_137;
  wire or_tmp_144;
  wire not_tmp_388;
  wire or_tmp_155;
  wire or_tmp_161;
  wire and_dcpl_674;
  wire or_tmp_175;
  wire or_tmp_177;
  wire mux_tmp_160;
  wire not_tmp_393;
  wire or_tmp_182;
  wire or_tmp_187;
  wire or_tmp_190;
  wire mux_tmp_171;
  wire or_tmp_194;
  wire or_tmp_200;
  wire or_tmp_206;
  wire and_dcpl_677;
  wire nor_tmp_116;
  wire mux_tmp_192;
  wire and_dcpl_678;
  wire and_dcpl_680;
  wire and_dcpl_681;
  wire and_dcpl_684;
  wire mux_tmp_195;
  wire and_dcpl_686;
  wire and_dcpl_689;
  wire and_dcpl_690;
  wire and_dcpl_693;
  wire and_dcpl_695;
  wire nor_tmp_121;
  wire or_tmp_228;
  wire or_tmp_229;
  wire or_tmp_230;
  wire nor_tmp_125;
  wire or_tmp_231;
  wire or_tmp_232;
  wire mux_tmp_199;
  wire and_dcpl_696;
  wire and_dcpl_697;
  wire mux_tmp_202;
  wire and_dcpl_703;
  wire nor_tmp_127;
  wire or_tmp_245;
  wire or_tmp_247;
  wire or_tmp_250;
  wire mux_tmp_215;
  wire or_tmp_259;
  wire or_tmp_267;
  wire or_tmp_268;
  wire or_tmp_269;
  wire or_tmp_272;
  wire or_tmp_273;
  wire mux_tmp_234;
  wire or_tmp_284;
  wire mux_tmp_244;
  wire or_tmp_291;
  wire and_dcpl_705;
  wire or_tmp_304;
  wire mux_tmp_255;
  wire and_dcpl_707;
  wire and_dcpl_710;
  wire and_dcpl_711;
  wire and_dcpl_714;
  wire and_dcpl_718;
  wire and_dcpl_719;
  wire and_dcpl_722;
  wire or_dcpl_308;
  wire [3:0] pe_config_manager_counter_sva_mx1;
  wire [4:0] operator_4_false_acc_sdt_sva_1;
  wire [5:0] nl_operator_4_false_acc_sdt_sva_1;
  reg [3:0] pe_config_num_manager_sva;
  wire state_0_sva_mx1;
  wire while_if_and_tmp_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiWrite_switch_lp_nor_tmp_1;
  reg pe_config_is_valid_sva;
  reg pe_config_is_zero_first_sva;
  reg pe_manager_zero_active_sva;
  reg pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  reg pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  reg PECore_UpdateFSM_switch_lp_and_7_itm_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
  reg PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  reg [8:0] operator_8_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_8_false_acc_sdt_sva_1;
  wire PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  wire PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1;
  reg PECore_RunFSM_switch_lp_nor_tmp_1;
  reg [1:0] state_2_1_sva;
  reg state_0_sva;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0;
  reg PECore_RunFSM_switch_lp_equal_tmp_1_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2;
  reg weight_mem_run_3_for_land_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg input_read_req_valid_lpi_1_dfm_1_10;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8;
  reg rva_in_reg_rw_sva_10;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_10;
  wire PECore_RunScale_if_for_1_operator_32_true_slc_32_1_svs_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_10;
  wire PECore_RunScale_if_for_2_operator_32_true_slc_32_1_svs_1;
  wire PECore_RunScale_if_for_3_operator_32_true_slc_32_1_svs_1;
  wire PECore_RunScale_if_for_4_operator_32_true_slc_32_1_svs_1;
  wire PECore_RunScale_if_for_5_operator_32_true_slc_32_1_svs_1;
  wire PECore_RunScale_if_for_7_operator_32_true_slc_32_1_svs_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_10;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  wire PECore_UpdateFSM_switch_lp_equal_tmp_6;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  wire PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
  wire PECore_UpdateFSM_switch_lp_nor_tmp_1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
  wire [7:0] pe_config_input_counter_sva_mx1;
  wire [8:0] operator_16_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_16_false_acc_sdt_sva_1;
  reg [7:0] pe_manager_num_input_sva;
  reg [7:0] pe_config_num_output_sva;
  wire PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8;
  reg weight_mem_run_3_for_land_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  wire PECore_RunScale_if_for_6_operator_32_true_slc_32_1_svs_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_9;
  wire PECore_RunScale_if_for_8_operator_32_true_slc_32_1_svs_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_9;
  wire PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  reg PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
  wire weight_mem_run_3_for_land_lpi_1_dfm_1_1;
  wire weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  wire weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_145_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_164_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_133_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_5_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_4_itm_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
  wire weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_127_sva_1;
  reg input_write_req_valid_lpi_1_dfm_1_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1;
  wire input_write_req_valid_lpi_1_dfm_5;
  wire input_mem_banks_write_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1;
  reg [14:0] pe_manager_base_input_sva;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1;
  reg rva_in_reg_rw_sva_5;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_4;
  wire PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3;
  reg rva_in_reg_rw_sva_st_1_10;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10;
  reg while_stage_0_12;
  reg rva_in_reg_rw_sva_9;
  reg input_read_req_valid_lpi_1_dfm_1_9;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
  reg rva_in_reg_rw_sva_st_1_9;
  reg rva_in_reg_rw_sva_st_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
  reg while_stage_0_11;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_8;
  reg while_stage_0_10;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
  reg while_stage_0_9;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  reg rva_in_reg_rw_sva_st_1_6;
  reg rva_in_reg_rw_sva_st_1_5;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  reg while_stage_0_7;
  reg while_stage_0_6;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_1;
  reg while_stage_0_5;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3;
  reg while_stage_0_4;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0;
  reg while_stage_0_3;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1;
  reg PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_1;
  reg rva_in_reg_rw_sva_st_1_4;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52;
  reg rva_in_reg_rw_sva_st_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  reg input_read_req_valid_lpi_1_dfm_1_8;
  reg rva_in_reg_rw_sva_st_1_8;
  reg rva_in_reg_rw_sva_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1;
  reg rva_in_reg_rw_sva_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg rva_in_reg_rw_sva_st_7;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  reg input_read_req_valid_lpi_1_dfm_1_7;
  reg rva_in_reg_rw_sva_st_1_7;
  reg rva_in_reg_rw_sva_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
  reg rva_in_reg_rw_sva_st_6;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
  reg input_read_req_valid_lpi_1_dfm_1_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
  reg while_stage_0_8;
  reg rva_in_reg_rw_sva_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
  reg rva_in_reg_rw_sva_st_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
  reg rva_in_reg_rw_sva_3;
  reg rva_in_reg_rw_sva_st_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
  reg rva_in_reg_rw_sva_st_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2;
  reg input_read_req_valid_lpi_1_dfm_1_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
  reg input_read_req_valid_lpi_1_dfm_1_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
  reg input_read_req_valid_lpi_1_dfm_1_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1;
  reg [3:0] while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9;
  reg weight_mem_run_3_for_5_and_28_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3;
  reg weight_mem_run_3_for_5_and_22_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5;
  reg [1:0] state_2_1_sva_dfm_1;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_2;
  reg while_and_1145_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_7_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  reg [7:0] weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_4_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_3_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_1_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_4_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs;
  wire operator_7_false_1_operator_7_false_1_or_mdf_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_3_2_0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_1_lpi_1_dfm_3_2_0;
  reg [14:0] weight_read_addrs_7_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_5_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_3_lpi_1_dfm_1;
  reg [2:0] weight_read_addrs_1_lpi_1_dfm_2_2_0;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  wire [11:0] nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  reg [14:0] pe_manager_base_weight_sva;
  reg [14:0] weight_read_addrs_1_lpi_1_dfm_1;
  wire [3:0] pe_manager_base_weight_sva_mx1_3_0;
  wire [14:0] pe_manager_base_weight_sva_mx2;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1;
  reg [7:0] while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4;
  wire [7:0] input_write_addrs_lpi_1_dfm_2;
  wire [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1;
  wire PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
  reg Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1;
  wire while_and_114_rgt;
  wire while_and_118_rgt;
  wire while_and_122_rgt;
  wire while_and_126_rgt;
  wire while_and_130_rgt;
  wire while_and_134_rgt;
  wire while_and_138_rgt;
  wire while_and_142_rgt;
  wire while_and_146_rgt;
  wire while_and_150_rgt;
  wire while_and_154_rgt;
  wire while_and_158_rgt;
  wire while_and_162_rgt;
  wire while_and_166_rgt;
  wire while_and_170_rgt;
  wire while_and_174_rgt;
  wire while_and_178_rgt;
  wire while_and_182_rgt;
  wire while_and_186_rgt;
  wire while_and_190_rgt;
  wire while_and_194_rgt;
  wire while_and_198_rgt;
  wire while_and_202_rgt;
  wire while_and_206_rgt;
  wire while_and_210_rgt;
  wire while_and_214_rgt;
  wire while_and_218_rgt;
  wire while_and_222_rgt;
  wire while_and_226_rgt;
  wire while_and_230_rgt;
  wire while_and_234_rgt;
  wire while_and_238_rgt;
  wire while_and_242_rgt;
  wire while_and_246_rgt;
  wire while_and_250_rgt;
  wire while_and_254_rgt;
  wire while_and_258_rgt;
  wire while_and_262_rgt;
  wire while_and_266_rgt;
  wire while_and_270_rgt;
  wire while_and_274_rgt;
  wire while_and_278_rgt;
  wire while_and_282_rgt;
  wire while_and_286_rgt;
  wire while_and_290_rgt;
  wire while_and_294_rgt;
  wire while_and_298_rgt;
  wire while_and_302_rgt;
  wire while_and_306_rgt;
  wire while_and_310_rgt;
  wire while_and_314_rgt;
  wire while_and_318_rgt;
  wire while_and_322_rgt;
  wire while_and_326_rgt;
  wire while_and_330_rgt;
  wire while_and_334_rgt;
  wire while_and_338_rgt;
  wire while_and_342_rgt;
  wire while_and_346_rgt;
  wire while_and_350_rgt;
  wire while_and_354_rgt;
  wire while_and_358_rgt;
  wire while_and_362_rgt;
  wire while_and_366_rgt;
  wire while_and_370_rgt;
  wire while_and_374_rgt;
  wire while_and_378_rgt;
  wire while_and_382_rgt;
  wire while_and_386_rgt;
  wire while_and_390_rgt;
  wire while_and_394_rgt;
  wire while_and_398_rgt;
  wire while_and_402_rgt;
  wire while_and_406_rgt;
  wire while_and_410_rgt;
  wire while_and_414_rgt;
  wire while_and_418_rgt;
  wire while_and_422_rgt;
  wire while_and_426_rgt;
  wire while_and_430_rgt;
  wire while_and_434_rgt;
  wire while_and_438_rgt;
  wire while_and_442_rgt;
  wire while_and_446_rgt;
  wire while_and_450_rgt;
  wire while_and_454_rgt;
  wire while_and_458_rgt;
  wire while_and_462_rgt;
  wire while_and_466_rgt;
  wire while_and_470_rgt;
  wire while_and_474_rgt;
  wire while_and_478_rgt;
  wire while_and_482_rgt;
  wire while_and_486_rgt;
  wire while_and_490_rgt;
  wire while_and_494_rgt;
  wire while_and_498_rgt;
  wire while_and_502_rgt;
  wire while_and_506_rgt;
  wire while_and_510_rgt;
  wire while_and_514_rgt;
  wire while_and_518_rgt;
  wire while_and_522_rgt;
  wire while_and_526_rgt;
  wire while_and_530_rgt;
  wire while_and_534_rgt;
  wire while_and_538_rgt;
  wire while_and_542_rgt;
  wire while_and_546_rgt;
  wire while_and_550_rgt;
  wire while_and_554_rgt;
  wire while_and_558_rgt;
  wire while_and_562_rgt;
  wire while_and_566_rgt;
  wire while_and_570_rgt;
  wire while_and_574_rgt;
  wire while_and_578_rgt;
  wire while_and_582_rgt;
  wire while_and_586_rgt;
  wire while_and_590_rgt;
  wire while_and_594_rgt;
  wire while_and_598_rgt;
  wire while_and_602_rgt;
  wire while_and_606_rgt;
  wire while_and_610_rgt;
  wire while_and_614_rgt;
  wire while_and_618_rgt;
  wire while_and_622_rgt;
  wire while_and_626_rgt;
  wire while_and_630_rgt;
  wire while_and_634_rgt;
  wire while_and_638_rgt;
  wire while_and_642_rgt;
  wire while_and_646_rgt;
  wire while_and_650_rgt;
  wire while_and_654_rgt;
  wire while_and_658_rgt;
  wire while_and_662_rgt;
  wire while_and_666_rgt;
  wire while_and_670_rgt;
  wire while_and_674_rgt;
  wire while_and_678_rgt;
  wire while_and_682_rgt;
  wire while_and_686_rgt;
  wire while_and_690_rgt;
  wire while_and_694_rgt;
  wire while_and_698_rgt;
  wire while_and_702_rgt;
  wire while_and_706_rgt;
  wire while_and_710_rgt;
  wire while_and_714_rgt;
  wire while_and_718_rgt;
  wire while_and_722_rgt;
  wire while_and_726_rgt;
  wire while_and_730_rgt;
  wire while_and_734_rgt;
  wire while_and_738_rgt;
  wire while_and_742_rgt;
  wire while_and_746_rgt;
  wire while_and_750_rgt;
  wire while_and_754_rgt;
  wire while_and_758_rgt;
  wire while_and_762_rgt;
  wire while_and_766_rgt;
  wire while_and_770_rgt;
  wire while_and_774_rgt;
  wire while_and_778_rgt;
  wire while_and_782_rgt;
  wire while_and_786_rgt;
  wire while_and_790_rgt;
  wire while_and_794_rgt;
  wire while_and_798_rgt;
  wire while_and_802_rgt;
  wire while_and_806_rgt;
  wire while_and_810_rgt;
  wire while_and_814_rgt;
  wire while_and_818_rgt;
  wire while_and_822_rgt;
  wire while_and_826_rgt;
  wire while_and_830_rgt;
  wire while_and_834_rgt;
  wire while_and_838_rgt;
  wire while_and_842_rgt;
  wire while_and_846_rgt;
  wire while_and_850_rgt;
  wire while_and_854_rgt;
  wire while_and_858_rgt;
  wire while_and_862_rgt;
  wire while_and_866_rgt;
  wire while_and_870_rgt;
  wire while_and_874_rgt;
  wire while_and_878_rgt;
  wire while_and_882_rgt;
  wire while_and_886_rgt;
  wire while_and_890_rgt;
  wire while_and_894_rgt;
  wire while_and_898_rgt;
  wire while_and_902_rgt;
  wire while_and_906_rgt;
  wire while_and_910_rgt;
  wire while_and_914_rgt;
  wire while_and_918_rgt;
  wire while_and_922_rgt;
  wire while_and_926_rgt;
  wire while_and_930_rgt;
  wire while_and_934_rgt;
  wire while_and_938_rgt;
  wire while_and_942_rgt;
  wire while_and_946_rgt;
  wire while_and_950_rgt;
  wire while_and_954_rgt;
  wire while_and_958_rgt;
  wire while_and_962_rgt;
  wire while_and_966_rgt;
  wire while_and_970_rgt;
  wire while_and_974_rgt;
  wire while_and_978_rgt;
  wire while_and_982_rgt;
  wire while_and_986_rgt;
  wire while_and_990_rgt;
  wire while_and_994_rgt;
  wire while_and_998_rgt;
  wire while_and_1002_rgt;
  wire while_and_1006_rgt;
  wire while_and_1010_rgt;
  wire while_and_1014_rgt;
  wire while_and_1018_rgt;
  wire while_and_1022_rgt;
  wire while_and_1026_rgt;
  wire while_and_1030_rgt;
  wire while_and_1034_rgt;
  wire while_and_1038_rgt;
  wire while_and_1042_rgt;
  wire while_and_1046_rgt;
  wire while_and_1050_rgt;
  wire while_and_1054_rgt;
  wire while_and_1058_rgt;
  wire while_and_1062_rgt;
  wire while_and_1066_rgt;
  wire while_and_1070_rgt;
  wire while_and_1074_rgt;
  wire while_and_1078_rgt;
  wire while_and_1082_rgt;
  wire while_and_1086_rgt;
  wire while_and_1090_rgt;
  wire while_and_1094_rgt;
  wire while_and_1098_rgt;
  wire while_and_1102_rgt;
  wire while_and_1106_rgt;
  wire while_and_1110_rgt;
  wire while_and_1114_rgt;
  wire while_and_1118_rgt;
  wire while_and_1122_rgt;
  wire while_and_1126_rgt;
  wire while_and_1130_rgt;
  wire while_and_1134_rgt;
  wire weight_mem_banks_read_1_for_mux_cse;
  wire weight_mem_banks_read_1_for_mux_1_cse;
  wire weight_mem_banks_read_1_for_mux_4_cse;
  wire weight_mem_banks_read_1_for_mux_5_cse;
  wire weight_mem_banks_read_1_for_mux_8_cse;
  wire weight_mem_banks_read_1_for_mux_9_cse;
  wire weight_mem_banks_read_1_for_mux_12_cse;
  wire weight_mem_banks_read_1_for_mux_13_cse;
  wire weight_mem_banks_read_1_for_mux_16_cse;
  wire weight_mem_banks_read_1_for_mux_17_cse;
  wire weight_mem_banks_read_1_for_mux_20_cse;
  wire weight_mem_banks_read_1_for_mux_21_cse;
  wire weight_mem_banks_read_1_for_mux_24_cse;
  wire weight_mem_banks_read_1_for_mux_25_cse;
  wire weight_mem_banks_read_1_for_mux_28_cse;
  wire weight_mem_banks_read_1_for_mux_29_cse;
  wire weight_mem_banks_write_if_for_if_mux_8_cse;
  wire weight_mem_banks_write_if_for_if_mux_9_cse;
  wire weight_mem_banks_read_for_mux_cse;
  wire weight_mem_banks_read_for_mux_1_cse;
  wire weight_mem_banks_write_if_for_if_mux_12_cse;
  wire weight_mem_banks_write_if_for_if_mux_13_cse;
  wire weight_mem_banks_read_for_mux_4_cse;
  wire weight_mem_banks_read_for_mux_5_cse;
  wire weight_mem_banks_write_if_for_if_mux_16_cse;
  wire weight_mem_banks_write_if_for_if_mux_17_cse;
  wire weight_mem_banks_read_for_mux_8_cse;
  wire weight_mem_banks_read_for_mux_9_cse;
  wire weight_mem_banks_write_if_for_if_mux_20_cse;
  wire weight_mem_banks_write_if_for_if_mux_21_cse;
  wire weight_mem_banks_read_for_mux_12_cse;
  wire weight_mem_banks_read_for_mux_13_cse;
  wire weight_mem_banks_write_if_for_if_mux_24_cse;
  wire weight_mem_banks_write_if_for_if_mux_25_cse;
  wire weight_mem_banks_read_for_mux_16_cse;
  wire weight_mem_banks_read_for_mux_17_cse;
  wire weight_mem_banks_write_if_for_if_mux_28_cse;
  wire weight_mem_banks_write_if_for_if_mux_29_cse;
  wire weight_mem_banks_read_for_mux_20_cse;
  wire weight_mem_banks_read_for_mux_21_cse;
  wire weight_mem_banks_write_if_for_if_mux_32_cse;
  wire weight_mem_banks_write_if_for_if_mux_33_cse;
  wire weight_mem_banks_read_for_mux_24_cse;
  wire weight_mem_banks_read_for_mux_25_cse;
  wire weight_mem_banks_write_if_for_if_mux_36_cse;
  wire weight_mem_banks_write_if_for_if_mux_37_cse;
  wire weight_mem_banks_read_for_mux_28_cse;
  wire weight_mem_banks_read_for_mux_29_cse;
  wire input_mem_banks_write_1_if_for_if_mux_cse;
  wire input_mem_banks_write_1_if_for_if_mux_1_cse;
  wire input_mem_banks_read_1_for_mux_cse;
  wire input_mem_banks_read_1_for_mux_1_cse;
  wire input_mem_banks_write_if_for_if_mux_cse;
  wire input_mem_banks_write_if_for_if_mux_1_cse;
  wire input_mem_banks_read_for_mux_cse;
  wire input_mem_banks_read_for_mux_1_cse;
  reg reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_31_cse;
  reg reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_30_cse;
  reg reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_7_cse;
  reg reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_3_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_act_port_Push_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire rva_out_reg_data_and_cse;
  wire accum_vector_data_and_cse;
  wire weight_port_read_out_data_and_1_cse;
  reg reg_rva_in_reg_rw_sva_st_1_1_cse;
  wire weight_port_read_out_data_and_28_cse;
  wire weight_port_read_out_data_and_32_cse;
  wire weight_port_read_out_data_and_40_cse;
  wire weight_port_read_out_data_and_48_cse;
  wire operator_15_false_1_and_cse;
  wire pe_config_num_manager_and_cse;
  wire PECore_DecodeAxiWrite_switch_lp_and_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
  wire or_202_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_cse;
  wire or_260_cse;
  wire or_253_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
  wire pe_manager_num_input_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_or_1_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_22_cse;
  wire Arbiter_8U_Roundrobin_pick_and_21_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_10_cse;
  wire Arbiter_8U_Roundrobin_pick_and_15_cse;
  wire [1:0] state_mux_1_cse;
  wire and_289_cse;
  wire and_562_cse;
  wire and_567_cse;
  wire PECore_RunMac_or_cse;
  wire and_741_cse;
  wire and_742_cse;
  wire and_740_cse;
  wire and_628_cse;
  wire and_733_cse;
  wire and_734_cse;
  wire or_111_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse;
  wire and_739_cse;
  wire and_751_cse;
  wire while_and_29_cse;
  wire nor_cse;
  wire nor_197_cse;
  wire nor_198_cse;
  wire nor_199_cse;
  wire nor_200_cse;
  wire nor_204_cse;
  wire nor_208_cse;
  wire and_129_cse;
  wire nor_218_cse;
  wire nor_219_cse;
  wire nor_216_cse;
  wire nor_217_cse;
  wire nand_17_cse;
  wire nor_275_cse;
  wire and_882_cse;
  wire and_881_cse;
  wire and_880_cse;
  wire and_886_cse;
  wire and_885_cse;
  wire and_884_cse;
  wire and_883_cse;
  wire and_887_cse;
  wire and_888_cse;
  wire and_893_cse;
  wire and_891_cse;
  wire and_890_cse;
  wire and_889_cse;
  wire and_896_cse;
  wire and_895_cse;
  wire and_894_cse;
  wire and_782_cse;
  wire and_897_cse;
  wire and_892_cse;
  wire and_812_cse;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_cse;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse;
  wire and_903_cse;
  wire and_910_cse;
  wire and_904_cse;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_cse;
  wire and_899_cse;
  wire and_901_cse;
  wire and_900_cse;
  wire and_898_cse;
  wire and_906_cse;
  wire and_908_cse;
  wire and_907_cse;
  wire and_905_cse;
  wire and_902_cse;
  wire and_909_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse;
  reg Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1;
  wire while_if_and_2_m1c;
  wire weight_mem_run_3_for_5_and_177_cse;
  wire pe_config_is_valid_and_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_cse;
  wire Arbiter_8U_Roundrobin_pick_and_23_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_35_cse;
  wire Arbiter_8U_Roundrobin_pick_and_35_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_46_cse;
  wire Arbiter_8U_Roundrobin_pick_and_43_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_58_cse;
  wire Arbiter_8U_Roundrobin_pick_and_49_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_70_cse;
  wire Arbiter_8U_Roundrobin_pick_and_55_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_82_cse;
  wire Arbiter_8U_Roundrobin_pick_and_61_cse;
  wire and_374_cse;
  wire pe_config_input_counter_and_cse;
  wire and_525_cse;
  wire and_108_cse;
  wire and_115_cse;
  wire and_122_cse;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1;
  wire PECore_DecodeAxiWrite_switch_lp_or_5_cse_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0;
  wire weight_mem_run_3_for_5_and_175_cse;
  wire weight_mem_run_3_for_5_and_176_cse;
  wire weight_mem_run_3_for_5_and_178_cse;
  wire weight_mem_run_3_for_5_and_179_cse;
  wire weight_mem_run_3_for_5_and_188_cse;
  wire weight_mem_run_3_for_5_and_181_cse;
  wire and_560_rmff;
  wire and_557_rmff;
  wire and_554_rmff;
  wire and_550_rmff;
  wire and_546_rmff;
  wire and_543_rmff;
  wire and_539_rmff;
  wire and_537_rmff;
  wire and_533_rmff;
  wire and_534_rmff;
  wire and_528_rmff;
  wire and_531_rmff;
  wire and_565_rmff;
  reg [34:0] accum_vector_data_0_34_0_sva;
  reg [34:0] accum_vector_data_7_34_0_sva;
  reg [34:0] accum_vector_data_6_34_0_sva;
  reg [34:0] accum_vector_data_5_34_0_sva;
  reg [34:0] accum_vector_data_4_34_0_sva;
  reg [34:0] accum_vector_data_3_34_0_sva;
  reg [34:0] accum_vector_data_2_34_0_sva;
  reg [34:0] accum_vector_data_1_34_0_sva;
  reg [7:0] pe_config_output_counter_sva;
  reg [7:0] pe_config_input_counter_sva;
  reg [31:0] act_port_reg_data_255_224_sva_dfm_1_1;
  wire [31:0] act_port_reg_data_223_192_sva_dfm_3;
  reg [31:0] act_port_reg_data_191_160_sva_dfm_1_1;
  wire [31:0] act_port_reg_data_159_128_sva_dfm_3;
  wire [31:0] act_port_reg_data_127_96_sva_dfm_3;
  wire [31:0] act_port_reg_data_95_64_sva_dfm_3;
  wire [31:0] act_port_reg_data_63_32_sva_dfm_3;
  wire [31:0] act_port_reg_data_31_0_sva_dfm_3;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_5;
  reg rva_out_reg_data_63_sva_dfm_4_5;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_5;
  reg rva_out_reg_data_47_sva_dfm_4_5;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_5;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_5;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_5;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_4;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0;
  reg weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
  reg [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1;
  reg [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1;
  reg [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1;
  reg weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
  wire [15:0] weight_port_read_out_data_7_1_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_7_0_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_7_3_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_7_2_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_7_5_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_7_4_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_7_7_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_7_6_sva_dfm_2;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_5;
  reg [15:0] weight_mem_run_3_for_5_mux_5_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_4_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_7_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_6_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_49_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_48_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_51_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_50_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_53_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_52_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_55_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_54_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_9_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_8_itm_1;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  reg [15:0] weight_port_read_out_data_1_7_sva_dfm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_14_itm_1;
  wire [15:0] weight_port_read_out_data_5_1_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_5_0_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_5_3_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_5_2_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_5_5_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_5_4_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_5_7_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_5_6_sva_dfm_2;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  reg [15:0] weight_port_read_out_data_2_1_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001;
  reg [15:0] weight_port_read_out_data_2_0_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002;
  reg [15:0] weight_port_read_out_data_2_3_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003;
  reg [15:0] weight_port_read_out_data_2_2_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000004;
  reg [15:0] weight_port_read_out_data_2_5_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000005;
  reg [15:0] weight_port_read_out_data_2_4_sva_dfm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_23_itm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000006;
  reg [15:0] weight_port_read_out_data_2_6_sva_dfm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_33_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_32_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_35_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_34_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_37_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_36_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_39_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_38_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_25_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_24_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_27_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_26_itm_1;
  reg [15:0] weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
  reg [14:0] weight_write_addrs_lpi_1_dfm_1_2;
  reg [15:0] weight_write_data_data_0_7_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_6_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_5_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_4_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_3_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_2_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_1_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_0_lpi_1_dfm_1_3_2;
  reg [11:0] weight_write_addrs_lpi_1_dfm_1_3_14_3;
  wire and_dcpl_723;
  wire or_dcpl;
  wire and_dcpl_724;
  wire mux_tmp_256;
  wire or_dcpl_309;
  wire nor_tmp_191;
  wire or_dcpl_314;
  wire or_dcpl_315;
  wire or_dcpl_316;
  wire and_647_ssc;
  wire and_648_ssc;
  wire and_649_ssc;
  reg [127:0] input_mem_banks_read_read_data_lpi_1_dfm_1_4;
  reg [127:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1;
  wire [127:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0;
  wire [111:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0;
  reg [1:0] weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_28;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_35;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1;
  wire or_639_tmp;
  wire mux_259_tmp;
  wire and_915_cse;
  wire and_916_cse;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_1_4;
  wire and_929_cse;
  wire and_930_cse;
  wire and_931_cse;
  wire and_932_cse;
  wire and_933_cse;
  wire and_934_cse;
  wire and_935_cse;
  wire nor_397_cse;
  wire and_947_cse;
  wire and_948_cse;
  wire and_949_cse;
  wire and_950_cse;
  wire and_951_cse;
  wire and_952_cse;
  wire nor_399_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55;
  wire mux_2_itm;
  wire mux_144_itm;
  wire mux_181_itm;
  wire mux_228_itm;
  wire mux_241_itm;
  reg weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_6_sva;
  reg [14:0] pe_manager_base_bias_sva;
  reg pe_config_is_cluster_sva;
  reg pe_config_is_bias_sva;
  reg [3:0] pe_config_manager_counter_sva;
  reg [31:0] act_port_reg_data_127_96_sva;
  reg [31:0] act_port_reg_data_159_128_sva;
  reg [31:0] act_port_reg_data_95_64_sva;
  reg [31:0] act_port_reg_data_191_160_sva;
  reg [31:0] act_port_reg_data_63_32_sva;
  reg [31:0] act_port_reg_data_223_192_sva;
  reg [31:0] act_port_reg_data_31_0_sva;
  reg [31:0] act_port_reg_data_255_224_sva;
  reg [15:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8;
  reg [127:0] input_mem_banks_bank_a_0_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_1_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_2_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_3_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_4_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_5_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_6_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_7_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_8_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_9_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_10_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_11_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_12_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_13_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_14_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_15_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_16_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_17_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_18_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_19_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_20_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_21_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_22_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_23_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_24_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_25_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_26_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_27_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_28_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_29_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_30_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_31_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_32_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_33_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_34_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_35_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_36_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_37_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_38_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_39_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_40_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_41_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_42_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_43_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_44_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_45_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_46_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_47_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_48_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_49_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_50_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_51_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_52_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_53_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_54_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_55_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_56_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_57_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_58_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_59_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_60_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_61_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_62_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_63_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_64_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_65_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_66_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_67_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_68_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_69_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_70_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_71_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_72_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_73_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_74_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_75_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_76_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_77_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_78_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_79_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_80_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_81_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_82_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_83_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_84_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_85_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_86_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_87_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_88_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_89_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_90_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_91_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_92_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_93_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_94_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_95_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_96_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_97_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_98_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_99_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_100_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_101_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_102_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_103_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_104_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_105_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_106_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_107_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_108_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_109_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_110_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_111_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_112_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_113_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_114_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_115_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_116_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_117_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_118_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_119_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_120_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_121_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_122_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_123_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_124_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_125_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_126_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_127_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_128_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_129_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_130_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_131_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_132_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_133_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_134_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_135_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_136_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_137_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_138_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_139_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_140_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_141_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_142_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_143_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_144_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_145_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_146_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_147_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_148_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_149_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_150_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_151_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_152_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_153_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_154_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_155_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_156_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_157_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_158_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_159_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_160_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_161_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_162_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_163_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_164_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_165_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_166_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_167_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_168_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_169_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_170_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_171_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_172_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_173_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_174_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_175_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_176_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_177_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_178_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_179_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_180_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_181_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_182_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_183_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_184_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_185_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_186_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_187_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_188_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_189_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_190_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_191_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_192_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_193_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_194_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_195_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_196_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_197_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_198_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_199_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_200_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_201_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_202_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_203_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_204_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_205_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_206_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_207_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_208_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_209_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_210_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_211_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_212_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_213_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_214_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_215_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_216_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_217_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_218_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_219_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_220_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_221_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_222_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_223_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_224_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_225_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_226_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_227_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_228_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_229_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_230_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_231_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_232_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_233_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_234_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_235_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_236_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_237_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_238_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_239_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_240_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_241_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_242_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_243_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_244_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_245_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_246_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_247_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_248_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_249_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_250_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_251_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_252_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_253_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_254_sva_dfm_2;
  reg [127:0] input_mem_banks_bank_a_255_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_4_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_5_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_6_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_7_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_1_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_2_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_4_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_4_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_4_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_4_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_4_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_4_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_4_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_4_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_7_sva_dfm_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_6;
  reg rva_out_reg_data_24_sva_dfm_6;
  reg rva_out_reg_data_31_sva_dfm_6;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_6;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_6;
  reg rva_out_reg_data_16_sva_dfm_6;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_6;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_6;
  reg rva_out_reg_data_8_sva_dfm_6;
  reg [6:0] rva_out_reg_data_7_1_sva_dfm_6;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_6;
  reg rva_out_reg_data_0_sva_dfm_6;
  reg [127:0] weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1;
  reg [127:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1;
  reg [127:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_6;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_6;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_6;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_6;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2;
  reg [3:0] pe_config_manager_counter_sva_dfm_3_1;
  reg [7:0] input_read_addrs_sva_1_1;
  wire [8:0] nl_input_read_addrs_sva_1_1;
  reg rva_out_reg_data_63_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_4;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_1;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_2;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_3;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_4;
  reg rva_out_reg_data_47_sva_dfm_4_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_3;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_4;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_1;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_2;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_3;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_4;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_1_2;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_5;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_5;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_5;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_1;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_2;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_4;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_5;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_6;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_7;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_8;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_9;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_10;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_1;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_2;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_3;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_4;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_5;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_6_1;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_7;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_8;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_2;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_3;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_4;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_5;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_6_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_7;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_8;
  reg [7:0] pe_config_output_counter_sva_dfm_1;
  reg [7:0] pe_config_input_counter_sva_dfm_1;
  reg [3:0] pe_config_manager_counter_sva_dfm_1;
  reg [127:0] rva_in_reg_data_sva_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
  reg [14:0] weight_write_addrs_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_0_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_1_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_2_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_3_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_4_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_5_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_6_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_7_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_2;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_1;
  reg [127:0] input_mem_banks_read_read_data_lpi_1_dfm_1_2;
  reg [127:0] input_mem_banks_read_read_data_lpi_1_dfm_1_3;
  reg [10:0] PEManager_15U_GetWeightAddr_else_acc_3_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
  reg [127:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  reg [14:0] pe_manager_base_weight_sva_dfm_3_1;
  reg [14:0] pe_manager_base_input_sva_dfm_3_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_36_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_37_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_39_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_31_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5;
  reg [15:0] weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1;
  reg [15:0] weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_1;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2;
  reg weight_mem_run_3_for_5_and_162_itm_1;
  reg weight_mem_run_3_for_5_and_163_itm_1;
  reg weight_mem_run_3_for_5_and_164_itm_1;
  reg weight_mem_run_3_for_5_and_164_itm_2;
  reg weight_mem_run_3_for_5_and_165_itm_1;
  reg weight_mem_run_3_for_5_and_166_itm_1;
  reg weight_mem_run_3_for_5_and_167_itm_1;
  reg weight_mem_run_3_for_5_and_168_itm_1;
  reg weight_mem_run_3_for_5_and_8_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
  reg weight_mem_run_3_for_5_and_15_itm_1;
  reg weight_mem_run_3_for_5_and_20_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1;
  reg weight_mem_run_3_for_5_and_30_itm_1;
  reg weight_mem_run_3_for_5_and_31_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_7_itm_1;
  reg weight_mem_run_3_for_5_and_60_itm_1;
  reg weight_mem_run_3_for_5_and_71_itm_1;
  reg weight_mem_run_3_for_5_and_86_itm_1;
  reg weight_mem_run_3_for_5_and_88_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2;
  reg weight_mem_run_3_for_5_and_92_itm_1;
  reg weight_mem_run_3_for_5_and_92_itm_2;
  reg weight_mem_run_3_for_5_and_94_itm_1;
  reg weight_mem_run_3_for_5_and_94_itm_2;
  reg weight_mem_run_3_for_5_and_95_itm_1;
  reg weight_mem_run_3_for_5_and_95_itm_2;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1;
  reg weight_mem_run_3_for_5_and_150_itm_1;
  reg weight_mem_run_3_for_5_and_150_itm_2;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_2;
  reg weight_mem_run_3_for_5_and_156_itm_1;
  reg weight_mem_run_3_for_5_and_156_itm_2;
  reg weight_mem_run_3_for_5_and_159_itm_1;
  reg weight_mem_run_3_for_5_and_159_itm_2;
  reg [34:0] ProductSum_for_acc_14_itm_1;
  wire [35:0] nl_ProductSum_for_acc_14_itm_1;
  reg [14:0] PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1;
  reg while_if_mux_19_itm_1;
  reg PECore_PushAxiRsp_mux_10_itm_1;
  reg PECore_PushAxiRsp_mux_18_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  reg [111:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_16;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_3_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0;
  wire [31:0] act_port_reg_data_255_224_sva_dfm_3;
  wire [31:0] act_port_reg_data_191_160_sva_dfm_3;
  wire PECore_PushAxiRsp_if_else_mux_18_mx0w2;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_mx0w0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_mx0w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0;
  wire weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0;
  wire weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0;
  wire weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
  wire [14:0] weight_read_addrs_1_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_3_lpi_1_dfm_1_1;
  wire [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_5_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_7_lpi_1_dfm_1_1;
  wire [3:0] pe_config_manager_counter_sva_mx0w0;
  wire [7:0] pe_config_output_counter_sva_mx1;
  wire pe_config_is_zero_first_sva_mx1;
  wire pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
  wire PECore_PushAxiRsp_if_else_mux_10_mx0w2;
  wire [15:0] rva_out_reg_data_127_112_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_111_96_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_95_80_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_79_64_sva_dfm_4_mx0w0;
  wire [14:0] rva_out_reg_data_62_48_sva_dfm_6_mx1;
  wire [6:0] rva_out_reg_data_46_40_sva_dfm_6_mx1;
  wire [3:0] rva_out_reg_data_39_36_sva_dfm_6_mx1;
  wire [3:0] rva_out_reg_data_35_32_sva_dfm_6_mx1;
  wire PECore_PushAxiRsp_mux_18_itm_1_mx0c1;
  wire [14:0] pe_manager_base_input_sva_mx1;
  wire PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  wire [15:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1;
  wire weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_mx0w0;
  wire nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_3_mux_mx0w1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_1;
  wire operator_3_false_1_operator_3_false_1_or_mdf_1_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1;
  wire operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_4;
  wire while_and_1148_cse_1;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000004;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000005;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000006;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_111_96_sva_1;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_95_80_sva_1;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_79_64_sva_1;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_63_48_sva_1;
  wire rva_out_reg_data_63_sva_dfm_7;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
  wire PECore_PushAxiRsp_if_asn_59;
  wire PECore_PushAxiRsp_if_asn_61;
  wire PECore_PushAxiRsp_if_asn_63;
  wire PECore_RunMac_asn_24;
  wire weight_mem_run_3_for_5_asn_290;
  wire weight_mem_run_3_for_5_asn_292;
  wire weight_mem_run_3_for_5_asn_294;
  wire weight_mem_run_3_for_5_asn_296;
  wire weight_mem_run_3_for_5_asn_298;
  wire weight_mem_run_3_for_5_asn_300;
  wire weight_mem_run_3_for_5_asn_302;
  wire weight_mem_run_3_for_5_asn_304;
  wire weight_mem_run_3_for_5_asn_306;
  wire weight_mem_run_3_for_5_asn_308;
  wire weight_mem_run_3_for_5_asn_310;
  wire weight_mem_run_3_for_5_asn_312;
  wire while_asn_631;
  wire PECore_PushAxiRsp_if_asn_67;
  wire PECore_PushAxiRsp_if_asn_69;
  wire PECore_PushAxiRsp_if_asn_71;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_96;
  wire weight_mem_run_3_for_5_and_166;
  wire weight_mem_run_3_for_5_and_168;
  wire weight_mem_run_3_for_5_and_172;
  wire weight_mem_run_3_for_5_and_174;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_57;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0;
  wire or_187_cse;
  wire PECore_PushAxiRsp_if_mux1h_9;
  wire [6:0] PECore_PushAxiRsp_if_mux1h_10;
  wire PECore_PushAxiRsp_if_mux1h_11;
  wire PECore_PushAxiRsp_if_mux1h_13;
  wire [6:0] PECore_PushAxiRsp_if_mux1h_14;
  wire PECore_PushAxiRsp_if_mux1h_15;
  wire [5:0] PECore_PushAxiRsp_if_mux1h_16;
  wire PECore_PushAxiRsp_if_mux1h_17;
  wire [15:0] weight_port_read_out_data_3_4_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_3_5_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_3_6_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_3_7_sva_dfm_3;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse;
  reg reg_rva_in_reg_rw_sva_2_cse;
  reg reg_weight_mem_run_3_for_5_and_20_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_15_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_30_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_162_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_163_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_165_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_166_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_168_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_167_itm_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse;
  wire weight_mem_banks_load_store_for_else_and_25_ssc;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_15;
  reg [14:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_14_0;
  wire weight_port_read_out_data_0_3_sva_dfm_mx0w3_15;
  wire [14:0] weight_port_read_out_data_0_3_sva_dfm_mx0w3_14_0;
  reg weight_port_read_out_data_0_1_sva_dfm_1_15;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_1_14_0;
  reg weight_port_read_out_data_0_1_sva_dfm_2_rsp_0;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_2_rsp_1;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd;
  reg [14:0] reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1;
  wire weight_port_read_out_data_0_1_sva_mx0_15;
  wire [14:0] weight_port_read_out_data_0_1_sva_mx0_14_0;
  wire and_654_ssc;
  wire and_656_ssc;
  wire and_657_ssc;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_15;
  reg [14:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_14_0;
  wire weight_mem_run_3_for_5_and_180_ssc;
  wire weight_port_read_out_data_and_64_ssc;
  reg weight_port_read_out_data_0_1_sva_dfm_1_1_15;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_1_1_14_0;
  reg weight_port_read_out_data_0_1_sva_15;
  reg [14:0] weight_port_read_out_data_0_1_sva_14_0;
  reg weight_port_read_out_data_0_1_sva_dfm_4_15;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_4_14_0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_ssc;
  wire weight_port_read_out_data_0_0_sva_dfm_mx0w1_15;
  wire [14:0] weight_port_read_out_data_0_0_sva_dfm_mx0w1_14_0;
  wire weight_port_read_out_data_0_3_sva_mx0_15;
  wire [14:0] weight_port_read_out_data_0_3_sva_mx0_14_0;
  wire and_964_ssc;
  wire weight_port_read_out_data_0_2_sva_dfm_mx0w1_15;
  wire [14:0] weight_port_read_out_data_0_2_sva_dfm_mx0w1_14_0;
  wire rva_out_reg_data_and_17_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_2_cse;
  wire rva_out_reg_data_and_20_cse;
  wire input_mem_banks_read_read_data_and_cse;
  wire weight_port_read_out_data_and_61_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_cse;
  wire act_port_reg_data_and_8_cse;
  wire PECore_PushOutput_if_and_cse;
  wire rva_in_reg_rw_and_cse;
  wire PECore_RunMac_if_and_1_cse;
  wire input_mem_banks_read_1_read_data_and_cse;
  wire weight_mem_run_3_for_aelse_and_cse;
  wire data_in_tmp_operator_2_for_and_1_cse;
  wire PECore_RunMac_if_and_5_cse;
  wire weight_mem_run_3_for_aelse_and_4_cse;
  wire weight_read_addrs_and_3_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_53_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_59_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_65_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_71_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_77_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_83_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_89_cse;
  wire weight_read_addrs_and_5_cse;
  wire weight_write_data_data_and_cse;
  wire weight_mem_write_arbxbar_xbar_for_1_for_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
  wire weight_read_addrs_and_7_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse;
  wire PECore_RunFSM_switch_lp_and_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_15_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_22_cse;
  wire Arbiter_8U_Roundrobin_pick_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_64_cse;
  wire weight_write_data_data_and_8_cse;
  wire rva_in_reg_rw_and_4_cse;
  wire PECore_UpdateFSM_switch_lp_and_11_cse;
  wire state_and_cse;
  wire weight_read_addrs_and_16_cse;
  wire weight_port_read_out_data_and_68_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_103_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_108_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_109_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse;
  wire weight_read_addrs_and_19_cse;
  wire while_if_and_11_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_24_cse;
  wire rva_in_reg_rw_and_6_cse;
  wire input_mem_banks_read_read_data_and_9_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse;
  wire while_if_and_15_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_7_cse;
  wire while_if_and_6_cse;
  wire rva_out_reg_data_and_30_cse;
  wire weight_port_read_out_data_and_72_cse;
  wire input_read_req_valid_and_1_cse;
  wire weight_mem_banks_load_store_for_else_and_cse;
  wire rva_in_reg_rw_and_2_cse;
  wire weight_mem_banks_load_store_for_else_and_24_cse;
  wire weight_mem_banks_load_store_for_else_and_27_cse;
  wire weight_mem_banks_load_store_for_else_and_28_cse;
  wire PECore_RunMac_if_and_2_cse;
  wire rva_in_reg_rw_and_9_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_117_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_122_cse;
  wire weight_read_addrs_and_24_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_83_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_89_cse;
  wire input_mem_banks_read_read_data_and_18_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse;
  wire pe_manager_base_weight_and_5_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_11_cse;
  wire while_if_and_7_cse;
  wire rva_out_reg_data_and_43_cse;
  wire weight_port_read_out_data_and_74_cse;
  wire input_read_req_valid_and_2_cse;
  wire PECore_UpdateFSM_switch_lp_and_10_cse;
  wire rva_in_reg_rw_and_5_cse;
  wire PECore_RunMac_if_and_3_cse;
  wire rva_in_reg_rw_and_12_cse;
  wire input_mem_banks_read_read_data_and_27_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_15_cse;
  wire while_if_and_8_cse;
  wire rva_out_reg_data_and_54_cse;
  wire input_read_req_valid_and_3_cse;
  wire PECore_UpdateFSM_switch_lp_and_17_cse;
  wire PECore_RunMac_if_and_4_cse;
  wire rva_in_reg_rw_and_15_cse;
  wire input_mem_banks_read_read_data_and_36_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_19_cse;
  wire rva_out_reg_data_and_65_cse;
  wire rva_out_reg_data_and_72_cse;
  wire PECore_UpdateFSM_switch_lp_and_18_cse;
  wire input_read_req_valid_and_4_cse;
  wire rva_out_reg_data_and_80_cse;
  wire PECore_RunMac_if_and_7_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_21_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_23_cse;
  wire rva_out_reg_data_and_87_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_27_cse;
  wire rva_out_reg_data_and_90_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse;
  wire rva_out_reg_data_and_97_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_35_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_36_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_40_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_45_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_49_cse;
  wire weight_port_read_out_data_and_76_cse;
  reg weight_port_read_out_data_0_1_sva_dfm_5_rsp_0;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_5_rsp_1;
  reg weight_port_read_out_data_0_3_sva_rsp_0;
  reg [14:0] weight_port_read_out_data_0_3_sva_rsp_1;
  wire weight_port_read_out_data_and_63_ssc;
  reg weight_port_read_out_data_0_0_sva_dfm_1_1_15;
  reg [14:0] weight_port_read_out_data_0_0_sva_dfm_1_1_14_0;
  wire weight_mem_run_3_for_5_and_195_ssc;
  reg weight_port_read_out_data_0_3_sva_dfm_1_1_15;
  reg [14:0] weight_port_read_out_data_0_3_sva_dfm_1_1_14_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_15;
  reg [14:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0;
  reg weight_port_read_out_data_0_0_sva_dfm_2_15;
  reg [14:0] weight_port_read_out_data_0_0_sva_dfm_2_14_0;
  reg weight_port_read_out_data_0_0_sva_dfm_2_15_1;
  reg [14:0] weight_port_read_out_data_0_0_sva_dfm_2_14_0_1;
  wire weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_15;
  wire [14:0] weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_14_0;
  wire weight_port_read_out_data_0_2_sva_mx0_15;
  wire [14:0] weight_port_read_out_data_0_2_sva_mx0_14_0;
  reg weight_port_read_out_data_0_2_sva_rsp_0;
  reg [14:0] weight_port_read_out_data_0_2_sva_rsp_1;
  reg weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
  reg [14:0] weight_port_read_out_data_0_0_sva_dfm_3_rsp_1;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_4_ftd;
  reg [14:0] reg_weight_port_read_out_data_0_0_sva_dfm_4_ftd_1;
  wire weight_mem_run_3_for_5_and_185_ssc;
  wire weight_mem_run_3_for_5_and_189_ssc;
  reg weight_port_read_out_data_0_2_sva_dfm_1_1_15;
  reg [14:0] weight_port_read_out_data_0_2_sva_dfm_1_1_14_0;
  reg weight_port_read_out_data_0_0_sva_dfm_5_15;
  reg [14:0] weight_port_read_out_data_0_0_sva_dfm_5_14_0;
  wire PECore_PushAxiRsp_if_mux1h_12_6;
  wire [5:0] PECore_PushAxiRsp_if_mux1h_12_5_0;
  reg rva_out_reg_data_15_9_sva_dfm_6_6;
  reg [5:0] rva_out_reg_data_15_9_sva_dfm_6_5_0;
  wire or_tmp_320;
  wire mux_tmp_268;
  wire not_tmp_469;
  wire or_dcpl_325;
  wire or_dcpl_336;
  wire or_dcpl_368;
  wire and_dcpl_891;
  wire or_tmp_374;
  wire or_tmp_406;
  wire or_tmp_407;
  wire mux_tmp_323;
  wire not_tmp_653;
  wire not_tmp_658;
  wire mux_tmp_335;
  wire not_tmp_662;
  wire or_tmp_425;
  wire and_tmp_24;
  wire or_647_cse;
  wire or_648_cse;
  wire or_649_cse;
  wire mux_289_cse;
  wire and_1066_cse;
  wire and_1090_cse;
  wire and_1085_cse;
  wire xor_5_cse;
  wire and_1118_cse;
  wire xor_13_cse;
  wire nor_431_cse;
  wire or_804_cse;
  wire and_1173_cse;
  wire and_1235_cse;
  wire and_1252_cse;
  wire and_1272_cse;
  wire nor_438_cse;
  wire nor_472_cse;
  wire and_1331_cse;
  wire nor_419_cse;
  wire nor_425_cse;
  wire nor_428_cse;
  wire nand_58_cse;
  wire or_691_cse;
  wire or_687_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse;
  wire and_1339_cse;
  wire and_985_cse;
  wire and_1053_cse;
  wire and_1179_cse;
  wire mux_347_cse;
  wire and_1062_cse;
  wire and_1086_cse;
  reg reg_rva_out_reg_data_15_9_sva_dfm_9_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_7_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_7_enexo;
  reg reg_rva_out_reg_data_127_112_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_111_96_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_95_80_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_4_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000001;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000002;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000003;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000004;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000005;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000006;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  reg reg_weight_read_addrs_6_14_1_lpi_1_dfm_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo;
  reg reg_weight_read_addrs_6_14_1_lpi_1_dfm_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1;
  reg reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_addrs_lpi_1_dfm_1_1_enexo;
  reg reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_config_num_output_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  reg reg_rva_in_reg_data_sva_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_127_112_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_111_96_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_95_80_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_4_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_127_112_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_111_96_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_95_80_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_4_2_enexo;
  reg reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_127_112_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_111_96_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_95_80_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_4_1_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_3;
  reg reg_rva_out_reg_data_30_25_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_4_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_1_3_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1;
  reg reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  reg reg_pe_manager_base_input_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_4_1_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_1_1_1_enexo;
  wire rva_out_reg_data_and_113_enex5;
  wire rva_out_reg_data_and_114_enex5;
  wire rva_out_reg_data_and_115_enex5;
  wire rva_out_reg_data_and_116_enex5;
  wire rva_out_reg_data_and_117_enex5;
  wire rva_out_reg_data_and_118_enex5;
  wire rva_out_reg_data_and_119_enex5;
  wire rva_out_reg_data_and_120_enex5;
  wire rva_out_reg_data_and_121_enex5;
  wire rva_out_reg_data_and_122_enex5;
  wire rva_out_reg_data_and_123_enex5;
  wire weight_port_read_out_data_and_78_enex5;
  wire input_mem_banks_read_read_data_and_48_enex5;
  wire input_mem_banks_read_read_data_and_49_enex5;
  wire input_mem_banks_read_read_data_and_50_enex5;
  wire input_mem_banks_read_read_data_and_51_enex5;
  wire input_mem_banks_read_1_read_data_and_5_enex5;
  wire weight_port_read_out_data_and_enex5;
  wire weight_port_read_out_data_and_79_enex5;
  wire weight_port_read_out_data_and_80_enex5;
  wire weight_port_read_out_data_and_81_enex5;
  wire weight_port_read_out_data_and_82_enex5;
  wire weight_port_read_out_data_and_83_enex5;
  wire weight_port_read_out_data_and_84_enex5;
  wire weight_port_read_out_data_and_85_enex5;
  wire input_mem_banks_read_1_read_data_and_1_enex5;
  wire weight_read_addrs_and_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5;
  wire weight_write_data_data_and_24_enex5;
  wire weight_write_data_data_and_25_enex5;
  wire weight_write_data_data_and_26_enex5;
  wire weight_write_data_data_and_27_enex5;
  wire weight_write_data_data_and_28_enex5;
  wire weight_write_data_data_and_29_enex5;
  wire weight_write_data_data_and_30_enex5;
  wire weight_write_data_data_and_31_enex5;
  wire weight_write_addrs_and_enex5;
  wire weight_write_data_data_and_32_enex5;
  wire weight_write_data_data_and_33_enex5;
  wire weight_write_data_data_and_34_enex5;
  wire weight_write_data_data_and_35_enex5;
  wire weight_write_data_data_and_36_enex5;
  wire weight_write_data_data_and_37_enex5;
  wire weight_write_data_data_and_38_enex5;
  wire weight_write_data_data_and_39_enex5;
  wire weight_write_addrs_and_3_enex5;
  wire weight_read_addrs_and_29_enex5;
  wire pe_config_UpdateManagerCounter_if_if_and_enex5;
  wire weight_read_addrs_and_30_enex5;
  wire PEManager_15U_PEManagerWrite_and_enex5;
  wire input_mem_banks_read_read_data_and_52_enex5;
  wire input_mem_banks_read_read_data_and_53_enex5;
  wire input_mem_banks_read_read_data_and_54_enex5;
  wire input_mem_banks_read_read_data_and_55_enex5;
  wire input_mem_banks_read_1_read_data_and_2_enex5;
  wire rva_out_reg_data_and_124_enex5;
  wire rva_out_reg_data_and_125_enex5;
  wire rva_out_reg_data_and_126_enex5;
  wire weight_port_read_out_data_and_86_enex5;
  wire rva_out_reg_data_and_127_enex5;
  wire rva_out_reg_data_and_128_enex5;
  wire rva_out_reg_data_and_129_enex5;
  wire rva_out_reg_data_and_130_enex5;
  wire rva_out_reg_data_and_131_enex5;
  wire rva_out_reg_data_and_132_enex5;
  wire rva_out_reg_data_and_133_enex5;
  wire rva_out_reg_data_and_134_enex5;
  wire input_mem_banks_read_read_data_and_56_enex5;
  wire input_mem_banks_read_read_data_and_57_enex5;
  wire input_mem_banks_read_read_data_and_58_enex5;
  wire input_mem_banks_read_read_data_and_59_enex5;
  wire input_mem_banks_read_1_read_data_and_3_enex5;
  wire rva_out_reg_data_and_135_enex5;
  wire rva_out_reg_data_and_136_enex5;
  wire rva_out_reg_data_and_137_enex5;
  wire weight_port_read_out_data_and_87_enex5;
  wire rva_out_reg_data_and_138_enex5;
  wire rva_out_reg_data_and_139_enex5;
  wire rva_out_reg_data_and_140_enex5;
  wire rva_out_reg_data_and_141_enex5;
  wire rva_out_reg_data_and_142_enex5;
  wire rva_out_reg_data_and_143_enex5;
  wire rva_out_reg_data_and_144_enex5;
  wire rva_out_reg_data_and_145_enex5;
  wire weight_mem_write_arbxbar_xbar_for_empty_and_enex5;
  wire input_mem_banks_read_read_data_and_60_enex5;
  wire input_mem_banks_read_read_data_and_61_enex5;
  wire input_mem_banks_read_read_data_and_62_enex5;
  wire input_mem_banks_read_read_data_and_63_enex5;
  wire rva_out_reg_data_and_146_enex5;
  wire rva_out_reg_data_and_147_enex5;
  wire rva_out_reg_data_and_148_enex5;
  wire rva_out_reg_data_and_149_enex5;
  wire rva_out_reg_data_and_150_enex5;
  wire rva_out_reg_data_and_151_enex5;
  wire rva_out_reg_data_and_152_enex5;
  wire rva_out_reg_data_and_153_enex5;
  wire rva_out_reg_data_and_154_enex5;
  wire rva_out_reg_data_and_155_enex5;
  wire rva_out_reg_data_and_156_enex5;
  wire input_mem_banks_read_read_data_and_64_enex5;
  wire input_mem_banks_read_read_data_and_65_enex5;
  wire input_mem_banks_read_read_data_and_66_enex5;
  wire input_mem_banks_read_read_data_and_67_enex5;
  wire rva_out_reg_data_and_157_enex5;
  wire rva_out_reg_data_and_158_enex5;
  wire rva_out_reg_data_and_159_enex5;
  wire rva_out_reg_data_and_160_enex5;
  wire rva_out_reg_data_and_161_enex5;
  wire rva_out_reg_data_and_162_enex5;
  wire rva_out_reg_data_and_163_enex5;
  wire rva_out_reg_data_and_164_enex5;
  wire rva_out_reg_data_and_165_enex5;
  wire input_mem_banks_read_read_data_and_46_enex5;
  wire rva_out_reg_data_and_166_enex5;
  wire rva_out_reg_data_and_167_enex5;
  wire rva_out_reg_data_and_168_enex5;
  wire rva_out_reg_data_and_169_enex5;
  wire rva_out_reg_data_and_170_enex5;
  wire rva_out_reg_data_and_171_enex5;
  wire rva_out_reg_data_and_172_enex5;
  wire input_mem_banks_read_read_data_and_47_enex5;
  wire rva_out_reg_data_and_173_enex5;
  wire rva_out_reg_data_and_174_enex5;
  wire rva_out_reg_data_and_175_enex5;
  wire rva_out_reg_data_and_176_enex5;
  wire rva_out_reg_data_and_177_enex5;
  wire rva_out_reg_data_and_104_enex5;
  wire rva_out_reg_data_and_178_enex5;
  wire rva_out_reg_data_and_179_enex5;
  wire rva_out_reg_data_and_180_enex5;
  wire rva_out_reg_data_and_181_enex5;
  wire weight_port_read_out_data_and_88_enex5;
  wire weight_port_read_out_data_and_89_enex5;
  wire weight_port_read_out_data_and_90_enex5;
  wire weight_port_read_out_data_and_91_enex5;
  wire weight_port_read_out_data_and_92_enex5;
  wire data_in_tmp_operator_2_for_and_tmp;
  wire rva_in_reg_data_and_tmp;
  wire input_mem_banks_read_1_read_data_and_4_tmp;
  wire input_mem_banks_read_read_data_and_45_tmp;
  wire pe_manager_base_input_and_tmp;
  wire and_1313_tmp;
  wire rva_in_reg_rw_and_3_cse;
  wire [34:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_1_itm;
  wire [34:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_2_itm;
  wire [34:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_3_itm;
  wire [34:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_4_itm;
  wire [34:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_5_itm;
  wire [34:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_6_itm;
  wire [34:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_7_itm;
  wire [34:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_itm;
  wire mux_335_itm;
  wire mux_256_cse;
  wire accum_vector_data_and_16_cse;
  wire accum_vector_data_and_17_cse;
  wire accum_vector_data_and_8_cse;
  wire accum_vector_data_and_14_cse;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27;
  wire mux_93_nl;
  wire and_877_nl;
  wire or_285_nl;
  wire mux_94_nl;
  wire nor_372_nl;
  wire or_289_nl;
  wire mux_98_nl;
  wire mux_97_nl;
  wire or_295_nl;
  wire or_293_nl;
  wire mux_95_nl;
  wire or_292_nl;
  wire or_291_nl;
  wire mux_101_nl;
  wire mux_100_nl;
  wire or_301_nl;
  wire or_300_nl;
  wire mux_105_nl;
  wire mux_104_nl;
  wire or_306_nl;
  wire or_305_nl;
  wire mux_108_nl;
  wire mux_107_nl;
  wire or_312_nl;
  wire or_311_nl;
  wire mux_111_nl;
  wire mux_110_nl;
  wire or_318_nl;
  wire or_636_nl;
  wire mux_114_nl;
  wire mux_113_nl;
  wire or_324_nl;
  wire or_323_nl;
  wire mux_117_nl;
  wire mux_116_nl;
  wire or_328_nl;
  wire or_327_nl;
  wire mux_121_nl;
  wire mux_120_nl;
  wire or_333_nl;
  wire or_332_nl;
  wire mux_128_nl;
  wire or_344_nl;
  wire mux_127_nl;
  wire and_564_nl;
  wire mux_126_nl;
  wire mux_125_nl;
  wire mux_124_nl;
  wire or_342_nl;
  wire mux_123_nl;
  wire or_341_nl;
  wire mux_122_nl;
  wire or_336_nl;
  wire mux_278_nl;
  wire and_984_nl;
  wire and_983_nl;
  wire PECore_UpdateFSM_switch_lp_not_27_nl;
  wire PECore_UpdateFSM_switch_lp_not_28_nl;
  wire PECore_UpdateFSM_switch_lp_not_29_nl;
  wire PECore_UpdateFSM_switch_lp_not_30_nl;
  wire PECore_UpdateFSM_switch_lp_not_31_nl;
  wire PECore_UpdateFSM_switch_lp_not_19_nl;
  wire mux_287_nl;
  wire mux_286_nl;
  wire mux_285_nl;
  wire[15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl;
  wire mux_288_nl;
  wire mux_301_nl;
  wire mux_300_nl;
  wire mux_307_nl;
  wire or_771_nl;
  wire mux_306_nl;
  wire mux_309_nl;
  wire mux_308_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_76_nl;
  wire mux_4_nl;
  wire nor_264_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_72_nl;
  wire mux_5_nl;
  wire nor_265_nl;
  wire mux_6_nl;
  wire or_22_nl;
  wire or_20_nl;
  wire mux_9_nl;
  wire mux_8_nl;
  wire or_27_nl;
  wire mux_7_nl;
  wire or_25_nl;
  wire or_23_nl;
  wire mux_10_nl;
  wire mux_311_nl;
  wire mux_310_nl;
  wire nor_429_nl;
  wire nor_430_nl;
  wire[10:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl;
  wire mux_31_nl;
  wire mux_30_nl;
  wire mux_29_nl;
  wire mux_28_nl;
  wire mux_17_nl;
  wire while_mux_1276_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl;
  wire mux_312_nl;
  wire[3:0] operator_4_false_acc_nl;
  wire[4:0] nl_operator_4_false_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_7_nl;
  wire mux_313_nl;
  wire mux_314_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_and_1_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_mux1h_15_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_nor_8_nl;
  wire mux_315_nl;
  wire and_1178_nl;
  wire and_1177_nl;
  wire or_814_nl;
  wire PECore_UpdateFSM_switch_lp_not_38_nl;
  wire PECore_UpdateFSM_switch_lp_not_21_nl;
  wire mux_3_nl;
  wire or_17_nl;
  wire or_16_nl;
  wire mux_35_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_2_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_20_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_24_nl;
  wire mux_36_nl;
  wire or_180_nl;
  wire mux_37_nl;
  wire or_181_nl;
  wire mux_38_nl;
  wire or_184_nl;
  wire mux_55_nl;
  wire or_201_nl;
  wire mux_54_nl;
  wire mux_53_nl;
  wire mux_52_nl;
  wire mux_51_nl;
  wire mux_50_nl;
  wire mux_49_nl;
  wire mux_48_nl;
  wire mux_47_nl;
  wire mux_46_nl;
  wire mux_373_nl;
  wire mux_45_nl;
  wire mux_43_nl;
  wire mux_39_nl;
  wire or_190_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_19_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_129_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_101_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_115_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_122_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_94_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_108_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_130_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_102_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_116_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_123_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_95_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_109_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_131_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_103_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_117_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_124_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_96_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_110_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_132_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_104_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_118_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_125_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_97_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_111_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_133_nl;
  wire[15:0] mux1h_2_nl;
  wire and_938_nl;
  wire and_939_nl;
  wire and_940_nl;
  wire not_1864_nl;
  wire mux_63_nl;
  wire mux_62_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_126_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_112_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl;
  wire or_641_nl;
  wire[15:0] mux_275_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_or_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_mux1h_37_nl;
  wire and_658_nl;
  wire and_660_nl;
  wire and_664_nl;
  wire and_668_nl;
  wire and_669_nl;
  wire and_661_nl;
  wire or_643_nl;
  wire nor_398_nl;
  wire mux_81_nl;
  wire mux_80_nl;
  wire mux_79_nl;
  wire mux_78_nl;
  wire mux_77_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_127_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_113_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_128_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_114_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_78_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_38_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_nl;
  wire mux_85_nl;
  wire[7:0] input_mem_banks_read_1_for_mux_nl;
  wire and_973_nl;
  wire mux_86_nl;
  wire weight_port_read_out_data_mux_18_nl;
  wire and_676_nl;
  wire nor_383_nl;
  wire mux_320_nl;
  wire mux_319_nl;
  wire mux_318_nl;
  wire mux_317_nl;
  wire or_868_nl;
  wire or_867_nl;
  wire or_866_nl;
  wire or_865_nl;
  wire or_864_nl;
  wire[14:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl;
  wire or_422_nl;
  wire weight_mem_run_3_for_5_and_158_nl;
  wire weight_mem_run_3_for_5_and_151_nl;
  wire weight_mem_run_3_for_5_and_100_nl;
  wire weight_mem_run_3_for_5_and_112_nl;
  wire mux_91_nl;
  wire nor_251_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl;
  wire PECore_RunScale_and_14_nl;
  wire PECore_RunScale_and_15_nl;
  wire PECore_RunScale_and_12_nl;
  wire PECore_RunScale_and_13_nl;
  wire PECore_RunScale_and_10_nl;
  wire PECore_RunScale_and_11_nl;
  wire PECore_RunScale_and_8_nl;
  wire PECore_RunScale_and_9_nl;
  wire PECore_RunScale_and_6_nl;
  wire PECore_RunScale_and_7_nl;
  wire PECore_RunScale_and_2_nl;
  wire PECore_RunScale_and_3_nl;
  wire weight_mem_run_3_for_5_and_36_nl;
  wire weight_mem_run_3_for_5_and_145_nl;
  wire PECore_RunScale_and_nl;
  wire PECore_RunScale_and_1_nl;
  wire PECore_RunScale_and_4_nl;
  wire PECore_RunScale_and_5_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_68_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_69_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_73_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_74_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_76_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_77_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_79_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_80_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_81_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_82_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_83_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_84_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_85_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_92_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_95_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_98_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_99_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_103_nl;
  wire[14:0] PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_nl;
  wire[14:0] nl_operator_15_false_acc_nl;
  wire[14:0] PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[12:0] operator_15_false_acc_1_nl;
  wire[13:0] nl_operator_15_false_acc_1_nl;
  wire[14:0] PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_2_nl;
  wire[14:0] nl_operator_15_false_acc_2_nl;
  wire[14:0] PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl;
  wire and_645_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl;
  wire and_638_nl;
  wire while_or_262_nl;
  wire while_and_2_nl;
  wire[7:0] pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl;
  wire[7:0] operator_8_false_acc_nl;
  wire[8:0] nl_operator_8_false_acc_nl;
  wire pe_config_UpdateInputCounter_not_nl;
  wire pe_config_input_counter_nand_nl;
  wire[7:0] pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl;
  wire[7:0] operator_8_false_1_acc_nl;
  wire[8:0] nl_operator_8_false_1_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_9_nl;
  wire pe_config_output_counter_nand_nl;
  wire while_and_75_nl;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl;
  wire while_if_or_nl;
  wire while_if_and_4_nl;
  wire PECore_PushAxiRsp_mux_24_nl;
  wire[15:0] while_if_while_if_and_16_nl;
  wire[15:0] while_if_while_if_and_17_nl;
  wire[15:0] while_if_while_if_and_18_nl;
  wire[15:0] while_if_while_if_and_19_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_nl;
  wire weight_mem_banks_load_store_1_for_else_else_or_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_4_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_6_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_8_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_2_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl;
  wire mux_159_nl;
  wire nor_384_nl;
  wire nor_385_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_6_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl;
  wire mux_189_nl;
  wire nor_386_nl;
  wire nor_387_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_24_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl;
  wire and_711_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_254_nl;
  wire or_613_nl;
  wire mux_253_nl;
  wire mux_252_nl;
  wire or_607_nl;
  wire mux_251_nl;
  wire or_595_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_44_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl;
  wire PECore_UpdateFSM_switch_lp_mux1h_14_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl;
  wire PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl;
  wire PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_89_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_81_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_73_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_87_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_80_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_88_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_81_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_89_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_82_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_90_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_83_nl;
  wire[7:0] PEManager_15U_GetInputAddr_acc_nl;
  wire[8:0] nl_PEManager_15U_GetInputAddr_acc_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_583_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_584_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_585_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_586_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_587_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_588_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_589_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_590_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_591_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_592_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_593_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_594_nl;
  wire or_11_nl;
  wire and_730_nl;
  wire or_103_nl;
  wire or_100_nl;
  wire or_110_nl;
  wire mux_26_nl;
  wire mux_25_nl;
  wire mux_24_nl;
  wire mux_23_nl;
  wire mux_22_nl;
  wire mux_21_nl;
  wire mux_20_nl;
  wire mux_372_nl;
  wire mux_19_nl;
  wire mux_34_nl;
  wire mux_33_nl;
  wire mux_32_nl;
  wire and_736_nl;
  wire or_205_nl;
  wire mux_64_nl;
  wire mux_66_nl;
  wire mux_74_nl;
  wire mux_73_nl;
  wire or_215_nl;
  wire or_213_nl;
  wire nor_285_nl;
  wire and_746_nl;
  wire nor_286_nl;
  wire or_304_nl;
  wire mux_103_nl;
  wire or_303_nl;
  wire mux_106_nl;
  wire or_308_nl;
  wire mux_109_nl;
  wire or_315_nl;
  wire mux_112_nl;
  wire or_320_nl;
  wire mux_115_nl;
  wire or_326_nl;
  wire or_331_nl;
  wire mux_119_nl;
  wire or_330_nl;
  wire mux_143_nl;
  wire mux_142_nl;
  wire mux_141_nl;
  wire nand_3_nl;
  wire mux_140_nl;
  wire mux_139_nl;
  wire mux_138_nl;
  wire nand_2_nl;
  wire nor_326_nl;
  wire mux_150_nl;
  wire mux_149_nl;
  wire mux_148_nl;
  wire or_435_nl;
  wire or_434_nl;
  wire nor_327_nl;
  wire mux_147_nl;
  wire mux_146_nl;
  wire mux_145_nl;
  wire or_428_nl;
  wire or_427_nl;
  wire mux_158_nl;
  wire mux_157_nl;
  wire mux_156_nl;
  wire mux_155_nl;
  wire nor_328_nl;
  wire nor_329_nl;
  wire nor_330_nl;
  wire nor_331_nl;
  wire mux_154_nl;
  wire mux_153_nl;
  wire mux_152_nl;
  wire nor_332_nl;
  wire nor_333_nl;
  wire nor_334_nl;
  wire nor_335_nl;
  wire or_463_nl;
  wire or_461_nl;
  wire nor_336_nl;
  wire mux_166_nl;
  wire mux_165_nl;
  wire mux_164_nl;
  wire nand_5_nl;
  wire nor_337_nl;
  wire mux_163_nl;
  wire mux_162_nl;
  wire mux_161_nl;
  wire nand_4_nl;
  wire mux_170_nl;
  wire mux_169_nl;
  wire mux_168_nl;
  wire or_470_nl;
  wire or_469_nl;
  wire or_468_nl;
  wire mux_174_nl;
  wire mux_173_nl;
  wire mux_172_nl;
  wire or_477_nl;
  wire or_476_nl;
  wire mux_180_nl;
  wire mux_179_nl;
  wire mux_178_nl;
  wire or_484_nl;
  wire or_483_nl;
  wire mux_177_nl;
  wire mux_176_nl;
  wire or_482_nl;
  wire or_481_nl;
  wire mux_175_nl;
  wire or_480_nl;
  wire or_473_nl;
  wire mux_188_nl;
  wire mux_187_nl;
  wire mux_186_nl;
  wire mux_185_nl;
  wire nor_338_nl;
  wire nor_339_nl;
  wire nor_340_nl;
  wire nor_341_nl;
  wire mux_184_nl;
  wire mux_183_nl;
  wire mux_182_nl;
  wire nor_342_nl;
  wire nor_343_nl;
  wire nor_344_nl;
  wire nor_345_nl;
  wire or_510_nl;
  wire mux_191_nl;
  wire or_509_nl;
  wire mux_190_nl;
  wire and_814_nl;
  wire or_508_nl;
  wire mux_194_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_605_nl;
  wire mux_198_nl;
  wire mux_197_nl;
  wire or_530_nl;
  wire mux_196_nl;
  wire or_524_nl;
  wire mux_201_nl;
  wire mux_200_nl;
  wire or_535_nl;
  wire or_534_nl;
  wire or_533_nl;
  wire or_532_nl;
  wire mux_208_nl;
  wire mux_207_nl;
  wire mux_206_nl;
  wire mux_205_nl;
  wire mux_204_nl;
  wire mux_203_nl;
  wire or_540_nl;
  wire or_539_nl;
  wire or_538_nl;
  wire or_537_nl;
  wire or_536_nl;
  wire mux_214_nl;
  wire mux_213_nl;
  wire mux_212_nl;
  wire or_550_nl;
  wire mux_211_nl;
  wire or_548_nl;
  wire mux_210_nl;
  wire mux_209_nl;
  wire or_546_nl;
  wire or_545_nl;
  wire or_543_nl;
  wire mux_218_nl;
  wire mux_217_nl;
  wire mux_216_nl;
  wire nand_7_nl;
  wire or_560_nl;
  wire mux_227_nl;
  wire mux_226_nl;
  wire mux_225_nl;
  wire nand_9_nl;
  wire mux_224_nl;
  wire mux_223_nl;
  wire or_558_nl;
  wire mux_222_nl;
  wire mux_221_nl;
  wire mux_220_nl;
  wire nand_8_nl;
  wire mux_219_nl;
  wire or_554_nl;
  wire mux_233_nl;
  wire or_577_nl;
  wire or_575_nl;
  wire mux_240_nl;
  wire mux_239_nl;
  wire mux_238_nl;
  wire mux_237_nl;
  wire mux_236_nl;
  wire or_580_nl;
  wire or_578_nl;
  wire mux_235_nl;
  wire or_574_nl;
  wire mux_232_nl;
  wire or_573_nl;
  wire or_572_nl;
  wire mux_231_nl;
  wire mux_230_nl;
  wire or_571_nl;
  wire mux_229_nl;
  wire or_561_nl;
  wire mux_243_nl;
  wire mux_242_nl;
  wire or_586_nl;
  wire or_585_nl;
  wire or_584_nl;
  wire or_583_nl;
  wire mux_250_nl;
  wire mux_249_nl;
  wire mux_248_nl;
  wire mux_247_nl;
  wire mux_246_nl;
  wire mux_245_nl;
  wire or_593_nl;
  wire or_592_nl;
  wire or_591_nl;
  wire or_590_nl;
  wire or_587_nl;
  wire while_mux_1335_nl;
  wire and_569_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl;
  wire weight_mem_banks_write_if_for_if_and_35_nl;
  wire weight_mem_banks_write_if_for_if_and_36_nl;
  wire weight_mem_banks_write_if_for_if_and_37_nl;
  wire weight_mem_banks_write_if_for_if_and_38_nl;
  wire weight_mem_banks_write_if_for_if_and_39_nl;
  wire weight_mem_banks_write_if_for_if_and_40_nl;
  wire weight_mem_banks_write_if_for_if_and_41_nl;
  wire weight_mem_banks_write_if_for_if_mux_7_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl;
  wire mux_136_nl;
  wire nor_381_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl;
  wire weight_mem_banks_write_if_for_if_and_28_nl;
  wire weight_mem_banks_write_if_for_if_and_29_nl;
  wire weight_mem_banks_write_if_for_if_and_30_nl;
  wire weight_mem_banks_write_if_for_if_and_31_nl;
  wire weight_mem_banks_write_if_for_if_and_32_nl;
  wire weight_mem_banks_write_if_for_if_and_33_nl;
  wire weight_mem_banks_write_if_for_if_and_34_nl;
  wire weight_mem_banks_write_if_for_if_mux_6_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl;
  wire mux_135_nl;
  wire nor_380_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl;
  wire weight_mem_banks_write_if_for_if_and_21_nl;
  wire weight_mem_banks_write_if_for_if_and_22_nl;
  wire weight_mem_banks_write_if_for_if_and_23_nl;
  wire weight_mem_banks_write_if_for_if_and_24_nl;
  wire weight_mem_banks_write_if_for_if_and_25_nl;
  wire weight_mem_banks_write_if_for_if_and_26_nl;
  wire weight_mem_banks_write_if_for_if_and_27_nl;
  wire weight_mem_banks_write_if_for_if_mux_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl;
  wire mux_134_nl;
  wire nor_379_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl;
  wire weight_mem_banks_write_if_for_if_and_14_nl;
  wire weight_mem_banks_write_if_for_if_and_15_nl;
  wire weight_mem_banks_write_if_for_if_and_16_nl;
  wire weight_mem_banks_write_if_for_if_and_17_nl;
  wire weight_mem_banks_write_if_for_if_and_18_nl;
  wire weight_mem_banks_write_if_for_if_and_19_nl;
  wire weight_mem_banks_write_if_for_if_and_20_nl;
  wire weight_mem_banks_write_if_for_if_mux_4_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl;
  wire mux_133_nl;
  wire nor_378_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl;
  wire weight_mem_banks_write_if_for_if_and_7_nl;
  wire weight_mem_banks_write_if_for_if_and_8_nl;
  wire weight_mem_banks_write_if_for_if_and_9_nl;
  wire weight_mem_banks_write_if_for_if_and_10_nl;
  wire weight_mem_banks_write_if_for_if_and_11_nl;
  wire weight_mem_banks_write_if_for_if_and_12_nl;
  wire weight_mem_banks_write_if_for_if_and_13_nl;
  wire weight_mem_banks_write_if_for_if_mux_3_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl;
  wire mux_132_nl;
  wire nor_377_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl;
  wire weight_mem_banks_write_if_for_if_and_nl;
  wire weight_mem_banks_write_if_for_if_and_1_nl;
  wire weight_mem_banks_write_if_for_if_and_2_nl;
  wire weight_mem_banks_write_if_for_if_and_3_nl;
  wire weight_mem_banks_write_if_for_if_and_4_nl;
  wire weight_mem_banks_write_if_for_if_and_5_nl;
  wire weight_mem_banks_write_if_for_if_and_6_nl;
  wire weight_mem_banks_write_if_for_if_mux_2_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl;
  wire mux_131_nl;
  wire nor_376_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_1_nl;
  wire weight_mem_banks_write_if_for_if_mux_54_nl;
  wire mux_130_nl;
  wire nor_375_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_nl;
  wire weight_mem_banks_write_if_for_if_mux_53_nl;
  wire mux_129_nl;
  wire nor_374_nl;
  wire PECore_PushAxiRsp_if_else_mux_19_nl;
  wire rva_out_reg_data_mux_25_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_21_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl;
  wire PECore_PushAxiRsp_if_else_mux_20_nl;
  wire rva_out_reg_data_mux_26_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_22_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_18_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_mux_25_nl;
  wire PECore_PushAxiRsp_if_else_mux_21_nl;
  wire rva_out_reg_data_mux_27_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_23_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_mux_19_nl;
  wire PECore_PushAxiRsp_if_else_mux_22_nl;
  wire rva_out_reg_data_mux_29_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_24_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_mux_20_nl;
  wire PECore_PushAxiRsp_if_else_mux_23_nl;
  wire rva_out_reg_data_mux_28_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl;
  wire[34:0] ProductSum_for_acc_25_nl;
  wire[35:0] nl_ProductSum_for_acc_25_nl;
  wire[34:0] ProductSum_for_acc_26_nl;
  wire[35:0] nl_ProductSum_for_acc_26_nl;
  wire[34:0] ProductSum_for_acc_27_nl;
  wire[35:0] nl_ProductSum_for_acc_27_nl;
  wire PECore_UpdateFSM_switch_lp_not_37_nl;
  wire[34:0] ProductSum_for_acc_19_nl;
  wire[35:0] nl_ProductSum_for_acc_19_nl;
  wire[34:0] ProductSum_for_acc_20_nl;
  wire[35:0] nl_ProductSum_for_acc_20_nl;
  wire[34:0] ProductSum_for_acc_21_nl;
  wire[35:0] nl_ProductSum_for_acc_21_nl;
  wire PECore_UpdateFSM_switch_lp_not_36_nl;
  wire[34:0] ProductSum_for_acc_13_nl;
  wire[35:0] nl_ProductSum_for_acc_13_nl;
  wire[34:0] ProductSum_for_acc_15_nl;
  wire[35:0] nl_ProductSum_for_acc_15_nl;
  wire PECore_UpdateFSM_switch_lp_not_35_nl;
  wire[34:0] ProductSum_for_acc_16_nl;
  wire[35:0] nl_ProductSum_for_acc_16_nl;
  wire[34:0] ProductSum_for_acc_17_nl;
  wire[35:0] nl_ProductSum_for_acc_17_nl;
  wire[34:0] ProductSum_for_acc_18_nl;
  wire[35:0] nl_ProductSum_for_acc_18_nl;
  wire PECore_UpdateFSM_switch_lp_not_34_nl;
  wire[34:0] ProductSum_for_acc_22_nl;
  wire[35:0] nl_ProductSum_for_acc_22_nl;
  wire[34:0] ProductSum_for_acc_23_nl;
  wire[35:0] nl_ProductSum_for_acc_23_nl;
  wire[34:0] ProductSum_for_acc_24_nl;
  wire[35:0] nl_ProductSum_for_acc_24_nl;
  wire PECore_UpdateFSM_switch_lp_not_23_nl;
  wire[34:0] ProductSum_for_acc_28_nl;
  wire[35:0] nl_ProductSum_for_acc_28_nl;
  wire[34:0] ProductSum_for_acc_29_nl;
  wire[35:0] nl_ProductSum_for_acc_29_nl;
  wire[34:0] ProductSum_for_acc_30_nl;
  wire[35:0] nl_ProductSum_for_acc_30_nl;
  wire PECore_UpdateFSM_switch_lp_not_33_nl;
  wire[34:0] ProductSum_for_acc_nl;
  wire[35:0] nl_ProductSum_for_acc_nl;
  wire[34:0] ProductSum_for_acc_34_nl;
  wire[35:0] nl_ProductSum_for_acc_34_nl;
  wire[34:0] ProductSum_for_acc_35_nl;
  wire[35:0] nl_ProductSum_for_acc_35_nl;
  wire PECore_UpdateFSM_switch_lp_not_39_nl;
  wire[34:0] ProductSum_for_acc_31_nl;
  wire[35:0] nl_ProductSum_for_acc_31_nl;
  wire[34:0] ProductSum_for_acc_32_nl;
  wire[35:0] nl_ProductSum_for_acc_32_nl;
  wire[34:0] ProductSum_for_acc_33_nl;
  wire[35:0] nl_ProductSum_for_acc_33_nl;
  wire PECore_UpdateFSM_switch_lp_not_32_nl;
  wire mux1h_1_nl;
  wire[14:0] mux1h_7_nl;
  wire not_1918_nl;
  wire mux_61_nl;
  wire mux_60_nl;
  wire mux_59_nl;
  wire mux_58_nl;
  wire mux_57_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_28_nl;
  wire[14:0] weight_mem_banks_load_store_for_else_mux1h_44_nl;
  wire not_1861_nl;
  wire mux1h_4_nl;
  wire[14:0] mux1h_6_nl;
  wire not_1917_nl;
  wire mux_342_nl;
  wire mux_341_nl;
  wire mux_340_nl;
  wire mux1h_3_nl;
  wire mux_72_nl;
  wire mux_71_nl;
  wire mux_70_nl;
  wire mux_69_nl;
  wire mux_68_nl;
  wire[14:0] mux1h_8_nl;
  wire not_1920_nl;
  wire mux_350_nl;
  wire mux_349_nl;
  wire or_903_nl;
  wire mux_348_nl;
  wire mux_344_nl;
  wire mux_343_nl;
  wire mux1h_nl;
  wire[14:0] mux1h_9_nl;
  wire not_1921_nl;
  wire mux1h_5_nl;
  wire[14:0] mux1h_10_nl;
  wire not_1923_nl;
  wire mux_1_nl;
  wire or_12_nl;
  wire mux_354_nl;
  wire mux_353_nl;
  wire mux_352_nl;
  wire mux_357_nl;
  wire or_916_nl;
  wire or_914_nl;
  wire mux_356_nl;
  wire mux_355_nl;
  wire and_1340_nl;
  wire and_1341_nl;
  wire and_1342_nl;
  wire weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl;
  wire mux_84_nl;
  wire mux_83_nl;
  wire mux_82_nl;
  wire[14:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_64_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_136_nl;
  wire mux_363_nl;
  wire mux_362_nl;
  wire nor_477_nl;
  wire mux_361_nl;
  wire or_688_nl;
  wire mux_334_nl;
  wire mux_333_nl;
  wire or_889_nl;
  wire or_888_nl;
  wire or_887_nl;
  wire or_892_nl;
  wire or_894_nl;
  wire nand_64_nl;
  wire or_901_nl;
  wire mux_346_nl;
  wire mux_345_nl;
  wire or_905_nl;
  wire mux_338_nl;
  wire mux_337_nl;
  wire and_1337_nl;
  wire mux_336_nl;
  wire and_1338_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [34:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_b = MUX_v_35_2_2(accum_vector_data_0_34_0_sva,
      PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_itm,
      accum_vector_data_and_16_cse);
  wire [34:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_b = MUX_v_35_2_2(accum_vector_data_7_34_0_sva,
      PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_7_itm,
      accum_vector_data_and_17_cse);
  wire [34:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_b = MUX_v_35_2_2(accum_vector_data_6_34_0_sva,
      PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_6_itm,
      accum_vector_data_and_16_cse);
  wire [34:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_b = MUX_v_35_2_2(accum_vector_data_5_34_0_sva,
      PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_5_itm,
      accum_vector_data_and_17_cse);
  wire [34:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_b = MUX_v_35_2_2(accum_vector_data_4_34_0_sva,
      PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_4_itm,
      accum_vector_data_and_16_cse);
  wire [34:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_b = MUX_v_35_2_2(accum_vector_data_3_34_0_sva,
      PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_3_itm,
      accum_vector_data_and_16_cse);
  wire [34:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_b = MUX_v_35_2_2(accum_vector_data_2_34_0_sva,
      PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_2_itm,
      accum_vector_data_and_16_cse);
  wire [34:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_b = MUX_v_35_2_2(accum_vector_data_1_34_0_sva,
      PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_1_itm,
      accum_vector_data_and_16_cse);
  wire  nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (~ reg_rva_in_reg_rw_sva_2_cse);
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0];
  wire  nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a = PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2
      & reg_rva_in_reg_rw_sva_2_cse;
  wire [2:0] nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s = weight_write_addrs_lpi_1_dfm_1_2[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s = {(weight_read_addrs_6_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_4[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s = weight_read_addrs_7_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s = {(weight_read_addrs_2_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s = {(weight_read_addrs_4_14_2_lpi_1_dfm_1_1[0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[1:0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s = weight_read_addrs_3_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s = weight_read_addrs_5_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s = weight_read_addrs_1_lpi_1_dfm_1_1[2:0];
  wire [255:0] nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun
      = {act_port_reg_data_255_224_sva_dfm_1_1 , act_port_reg_data_223_192_sva_dfm_3
      , act_port_reg_data_191_160_sva_dfm_1_1 , act_port_reg_data_159_128_sva_dfm_3
      , act_port_reg_data_127_96_sva_dfm_3 , act_port_reg_data_95_64_sva_dfm_3 ,
      act_port_reg_data_63_32_sva_dfm_3 , act_port_reg_data_31_0_sva_dfm_3};
  wire [127:0] nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun
      = {rva_out_reg_data_127_112_sva_dfm_4_5 , rva_out_reg_data_111_96_sva_dfm_4_5
      , rva_out_reg_data_95_80_sva_dfm_4_5 , rva_out_reg_data_79_64_sva_dfm_4_5 ,
      rva_out_reg_data_63_sva_dfm_4_5 , rva_out_reg_data_62_48_sva_dfm_4_5 , rva_out_reg_data_47_sva_dfm_4_5
      , rva_out_reg_data_46_40_sva_dfm_4_5 , rva_out_reg_data_39_36_sva_dfm_4_5 ,
      rva_out_reg_data_35_32_sva_dfm_4_5 , PECore_PushAxiRsp_if_mux1h_17 , PECore_PushAxiRsp_if_mux1h_16
      , PECore_PushAxiRsp_if_mux1h_15 , PECore_PushAxiRsp_if_mux1h_14 , PECore_PushAxiRsp_if_mux1h_13
      , PECore_PushAxiRsp_if_mux1h_12_6 , PECore_PushAxiRsp_if_mux1h_12_5_0 , PECore_PushAxiRsp_if_mux1h_11
      , PECore_PushAxiRsp_if_mux1h_10 , PECore_PushAxiRsp_if_mux1h_9};
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd35),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_b[34:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd35),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_b[34:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd35),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_b[34:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd35),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_b[34:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd35),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_b[34:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd35),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_b[34:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd35),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_b[34:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd35),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_b[34:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_z)
    );
  PECore_mgc_muladd1 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_cst(32'sd1),
  .signd_cst(32'sd0),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd11),
  .add_axb(32'sd1),
  .add_c(32'sd1),
  .add_d(32'sd1),
  .use_const(32'sd1)) PEManager_15U_GetWeightAddr_else_acc_4_cmp (
      .a(pe_config_output_counter_sva),
      .b(pe_manager_num_input_sva),
      .c(pe_config_input_counter_sva),
      .cst(1'b0),
      .z(PEManager_15U_GetWeightAddr_else_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_for_1_lshift_rg (
      .a(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a),
      .s(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_write_arbxbar_xbar_for_lshift_rg (
      .a(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a),
      .s(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s[2:0]),
      .z(weight_mem_write_arbxbar_xbar_for_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi PECore_PECoreRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(fsm_output)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi PECore_PECoreRun_input_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_oswt_pff(and_565_rmff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi PECore_PECoreRun_act_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(reg_act_port_Push_mioi_iswt0_cse),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun[255:0]),
      .act_port_Push_mioi_oswt_pff(and_567_cse)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi PECore_PECoreRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_oswt_pff(and_565_rmff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi PECore_PECoreRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun[127:0]),
      .rva_out_Push_mioi_oswt_pff(and_562_cse)
    );
  PECore_PECore_PECoreRun_wait_dp PECore_PECoreRun_wait_dp_inst (
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .PECoreRun_wen(PECoreRun_wen),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg(and_560_rmff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg(and_557_rmff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg(and_554_rmff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg(and_550_rmff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg(and_546_rmff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg(and_543_rmff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg(and_539_rmff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg(and_537_rmff),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo(reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_7_cse),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg(and_533_rmff),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_1(reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_3_cse),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg_1(and_534_rmff),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_cgo(reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_31_cse),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg(and_528_rmff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_5(reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_30_cse),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg_5(and_531_rmff)
    );
  PECore_PECore_PECoreRun_staller PECore_PECoreRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp)
    );
  PECore_PECore_PECoreRun_PECoreRun_fsm PECore_PECoreRun_PECoreRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .fsm_output(fsm_output)
    );
  assign weight_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_84);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign weight_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_84);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign weight_mem_banks_read_1_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_86);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign weight_mem_banks_read_1_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_86);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign weight_mem_banks_read_1_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_88);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 );
  assign weight_mem_banks_read_1_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_88);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign weight_mem_banks_read_1_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_90);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 );
  assign weight_mem_banks_read_1_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_90);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign weight_mem_banks_read_1_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_92);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 );
  assign weight_mem_banks_read_1_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_92);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign weight_mem_banks_read_1_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_94);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 );
  assign weight_mem_banks_read_1_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_94);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign weight_mem_banks_read_1_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_80);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 );
  assign weight_mem_banks_read_1_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_80);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign weight_mem_banks_read_1_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_82);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 );
  assign weight_mem_banks_read_1_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_82);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign weight_mem_banks_write_if_for_if_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_167);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 );
  assign weight_mem_banks_write_if_for_if_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_167);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign weight_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_168);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 );
  assign weight_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_168);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign weight_mem_banks_write_if_for_if_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_169);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 );
  assign weight_mem_banks_write_if_for_if_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_169);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1
      = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1
      = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign weight_mem_banks_read_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_170);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 );
  assign weight_mem_banks_read_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_170);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign weight_mem_banks_write_if_for_if_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_172);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 );
  assign weight_mem_banks_write_if_for_if_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_172);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2
      = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2
      = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign weight_mem_banks_read_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_173);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 );
  assign weight_mem_banks_read_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_173);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign weight_mem_banks_write_if_for_if_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_175);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 );
  assign weight_mem_banks_write_if_for_if_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_175);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3
      = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3
      = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign weight_mem_banks_read_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_176);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 );
  assign weight_mem_banks_read_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_176);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign weight_mem_banks_write_if_for_if_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_177);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 );
  assign weight_mem_banks_write_if_for_if_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_177);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4
      = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4
      = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign weight_mem_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_178);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 );
  assign weight_mem_banks_read_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_178);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign weight_mem_banks_write_if_for_if_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_179);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 );
  assign weight_mem_banks_write_if_for_if_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_179);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5
      = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5
      = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign weight_mem_banks_read_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_180);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 );
  assign weight_mem_banks_read_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_180);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign weight_mem_banks_write_if_for_if_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_182);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 );
  assign weight_mem_banks_write_if_for_if_mux_33_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_182);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6
      = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6
      = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign weight_mem_banks_read_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_183);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 );
  assign weight_mem_banks_read_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_183);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign weight_mem_banks_write_if_for_if_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_185);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 );
  assign weight_mem_banks_write_if_for_if_mux_37_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_185);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7
      = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7
      = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign weight_mem_banks_read_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_186);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 );
  assign weight_mem_banks_read_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_186);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign input_mem_banks_write_1_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_196);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 );
  assign input_mem_banks_write_1_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_196);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8
      = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_3 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8
      = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign input_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_193);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 );
  assign input_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_193);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign input_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_207);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 );
  assign input_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_207);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9
      = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_1 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9
      = input_mem_banks_write_if_for_if_mux_1_cse;
  assign input_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_210);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 );
  assign input_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_210);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign and_525_cse = and_dcpl_48 & PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  assign and_528_rmff = (and_dcpl_527 | and_525_cse | and_dcpl_523) & fsm_output;
  assign and_531_rmff = ((and_dcpl_35 & PECore_RunMac_PECore_RunMac_if_and_svs_8)
      | and_dcpl_527 | and_dcpl_523) & fsm_output;
  assign and_877_nl = (~(while_stage_0_11 & PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9))
      & or_tmp_79;
  assign or_285_nl = PECore_RunMac_PECore_RunMac_if_and_svs_9 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9;
  assign mux_93_nl = MUX_s_1_2_2(and_877_nl, or_tmp_79, or_285_nl);
  assign and_533_rmff = (~ mux_93_nl) & fsm_output;
  assign nor_372_nl = ~(while_stage_0_9 | (~ or_tmp_79));
  assign or_289_nl = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7) | PECore_RunMac_PECore_RunMac_if_and_svs_st_7
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  assign mux_94_nl = MUX_s_1_2_2(nor_372_nl, or_tmp_79, or_289_nl);
  assign and_534_rmff = (~ mux_94_nl) & fsm_output;
  assign or_295_nl = weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | not_tmp_249;
  assign or_292_nl = nor_tmp_17 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_1;
  assign or_291_nl = (~(weight_mem_run_3_for_5_and_28_itm_1 | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3)
      | (~ while_stage_0_7))) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_1;
  assign mux_95_nl = MUX_s_1_2_2(or_292_nl, or_291_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_293_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
      | mux_95_nl;
  assign mux_97_nl = MUX_s_1_2_2(or_295_nl, or_293_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_98_nl = MUX_s_1_2_2(not_tmp_249, mux_97_nl, while_stage_0_6);
  assign and_537_rmff = (mux_98_nl | and_dcpl_536) & fsm_output;
  assign or_301_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | not_tmp_252;
  assign or_300_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 | not_tmp_252;
  assign mux_100_nl = MUX_s_1_2_2(or_301_nl, or_300_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_101_nl = MUX_s_1_2_2(not_tmp_252, mux_100_nl, while_stage_0_6);
  assign and_539_rmff = (mux_101_nl | and_dcpl_538) & fsm_output;
  assign or_306_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp;
  assign or_305_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2)))
      | and_tmp;
  assign mux_104_nl = MUX_s_1_2_2(or_306_nl, or_305_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_105_nl = MUX_s_1_2_2(and_tmp, mux_104_nl, while_stage_0_6);
  assign and_543_rmff = (mux_105_nl | and_dcpl_179) & fsm_output;
  assign or_312_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_1;
  assign or_311_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2)))
      | and_tmp_1;
  assign mux_107_nl = MUX_s_1_2_2(or_312_nl, or_311_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_108_nl = MUX_s_1_2_2(and_tmp_1, mux_107_nl, while_stage_0_6);
  assign and_546_rmff = (mux_108_nl | and_dcpl_177) & fsm_output;
  assign or_318_nl = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_2;
  assign or_636_nl = (~((~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1)) | and_tmp_2;
  assign mux_110_nl = MUX_s_1_2_2(or_318_nl, or_636_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_111_nl = MUX_s_1_2_2(and_tmp_2, mux_110_nl, while_stage_0_6);
  assign and_550_rmff = (mux_111_nl | and_dcpl_175) & fsm_output;
  assign or_324_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_3;
  assign or_323_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse)))
      | and_tmp_3;
  assign mux_113_nl = MUX_s_1_2_2(or_324_nl, or_323_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_114_nl = MUX_s_1_2_2(and_tmp_3, mux_113_nl, while_stage_0_6);
  assign and_554_rmff = (mux_114_nl | and_dcpl_172) & fsm_output;
  assign or_328_nl = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_4;
  assign or_327_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse)))
      | and_tmp_4;
  assign mux_116_nl = MUX_s_1_2_2(or_328_nl, or_327_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_117_nl = MUX_s_1_2_2(and_tmp_4, mux_116_nl, while_stage_0_6);
  assign and_557_rmff = (mux_117_nl | and_dcpl_169) & fsm_output;
  assign or_333_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_5;
  assign or_332_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse)))
      | and_tmp_5;
  assign mux_120_nl = MUX_s_1_2_2(or_333_nl, or_332_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_121_nl = MUX_s_1_2_2(and_tmp_5, mux_120_nl, while_stage_0_6);
  assign and_560_rmff = (mux_121_nl | and_dcpl_167) & fsm_output;
  assign or_342_nl = (start_PopNB_mioi_data_rsc_z_mxwt & start_PopNB_mioi_return_rsc_z_mxwt
      & pe_config_is_valid_sva & PECore_UpdateFSM_switch_lp_and_7_itm_1) | or_tmp_121;
  assign mux_124_nl = MUX_s_1_2_2(or_342_nl, or_tmp_123, state_2_1_sva[1]);
  assign or_341_nl = (~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1)
      | pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8])
      | or_tmp_123;
  assign mux_123_nl = MUX_s_1_2_2(nand_tmp_1, or_341_nl, state_2_1_sva[1]);
  assign mux_125_nl = MUX_s_1_2_2(mux_124_nl, mux_123_nl, PECore_UpdateFSM_switch_lp_equal_tmp_5_1);
  assign mux_122_nl = MUX_s_1_2_2(or_tmp_123, nand_tmp_1, PECore_UpdateFSM_switch_lp_equal_tmp_5_1);
  assign or_336_nl = state_0_sva | (state_2_1_sva[0]);
  assign mux_126_nl = MUX_s_1_2_2(mux_125_nl, mux_122_nl, or_336_nl);
  assign and_564_nl = PECore_UpdateFSM_switch_lp_nor_7_itm_1 & ((PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      & pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1)
      | mux_126_nl);
  assign mux_127_nl = MUX_s_1_2_2(and_564_nl, state_0_sva, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign or_344_nl = (state_2_1_sva_dfm_1!=2'b00) | mux_127_nl;
  assign mux_128_nl = MUX_s_1_2_2(or_tmp_129, or_344_nl, while_stage_0_3);
  assign and_565_rmff = (~ mux_128_nl) & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign PECore_DecodeAxiRead_switch_lp_and_2_cse = PECoreRun_wen & and_dcpl_7 &
      (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 | input_read_req_valid_lpi_1_dfm_1_9
      | rva_in_reg_rw_sva_9));
  assign rva_out_reg_data_and_17_cse = PECoreRun_wen & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_9
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9)) & while_stage_0_11 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9
      & (~ rva_in_reg_rw_sva_st_1_9) & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7)
      & and_dcpl_10 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9) & (~ rva_in_reg_rw_sva_st_9)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
  assign rva_out_reg_data_and_113_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_15_9_sva_dfm_9_enexo;
  assign rva_out_reg_data_and_114_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_23_17_sva_dfm_7_enexo;
  assign rva_out_reg_data_and_115_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_30_25_sva_dfm_7_enexo;
  assign rva_out_reg_data_and_20_cse = PECoreRun_wen & and_dcpl_7;
  assign rva_out_reg_data_and_116_enex5 = rva_out_reg_data_and_20_cse & reg_rva_out_reg_data_127_112_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_117_enex5 = rva_out_reg_data_and_20_cse & reg_rva_out_reg_data_111_96_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_118_enex5 = rva_out_reg_data_and_20_cse & reg_rva_out_reg_data_95_80_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_119_enex5 = rva_out_reg_data_and_20_cse & reg_rva_out_reg_data_79_64_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_120_enex5 = rva_out_reg_data_and_20_cse & reg_rva_out_reg_data_62_48_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_121_enex5 = rva_out_reg_data_and_20_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_122_enex5 = rva_out_reg_data_and_20_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_123_enex5 = rva_out_reg_data_and_20_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo;
  assign input_mem_banks_read_read_data_and_cse = PECoreRun_wen & and_dcpl_7 & (~
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7) & input_read_req_valid_lpi_1_dfm_1_9;
  assign weight_port_read_out_data_and_61_cse = PECoreRun_wen & and_dcpl_6 & (~ rva_in_reg_rw_sva_st_1_9)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
  assign weight_port_read_out_data_and_78_enex5 = weight_port_read_out_data_and_61_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_cse = PECoreRun_wen & (~((~(while_stage_0_12 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10))
      | rva_in_reg_rw_sva_10 | (~ fsm_output)));
  assign input_mem_banks_read_read_data_and_48_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo;
  assign input_mem_banks_read_read_data_and_49_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo;
  assign input_mem_banks_read_read_data_and_50_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo;
  assign input_mem_banks_read_read_data_and_51_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo;
  assign rva_in_reg_rw_and_cse = PECoreRun_wen & while_stage_0_11;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_cse = PECoreRun_wen & and_dcpl_6
      & (~(rva_in_reg_rw_sva_st_1_9 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7))
      & and_dcpl_10 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
  assign act_port_reg_data_and_8_cse = PECoreRun_wen & and_dcpl_28 & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  assign PECore_PushOutput_if_and_cse = PECoreRun_wen & and_dcpl_28;
  assign or_649_cse = (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9) | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  assign and_984_nl = ((~ while_stage_0_11) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9)
      & or_tmp_320;
  assign and_983_nl = ((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_9) | PECore_RunMac_PECore_RunMac_if_and_svs_9
      | (~ while_stage_0_11) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9)
      & or_tmp_320;
  assign mux_278_nl = MUX_s_1_2_2(and_984_nl, and_983_nl, or_649_cse);
  assign and_985_cse = mux_278_nl & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10)
      & while_stage_0_12 & PECoreRun_wen;
  assign accum_vector_data_and_cse = PECoreRun_wen & fsm_output;
  assign accum_vector_data_and_8_cse = or_647_cse & while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9)
      & fsm_output & PECoreRun_wen & (~ or_dcpl_314);
  assign PECore_RunMac_if_and_1_cse = PECoreRun_wen & and_dcpl_35;
  assign while_if_and_6_cse = PECoreRun_wen & while_stage_0_10;
  assign accum_vector_data_and_14_cse = or_648_cse & while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8)
      & fsm_output & PECoreRun_wen & (~ or_dcpl_315);
  assign PECore_RunMac_if_and_2_cse = PECoreRun_wen & (and_dcpl_41 | and_dcpl_325);
  assign PECore_UpdateFSM_switch_lp_and_10_cse = PECoreRun_wen & and_dcpl_41;
  assign while_if_and_7_cse = PECoreRun_wen & while_stage_0_9;
  assign PECore_RunMac_if_and_3_cse = PECoreRun_wen & (~(rva_in_reg_rw_sva_st_1_6
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6))
      & while_stage_0_8;
  assign while_if_and_8_cse = PECoreRun_wen & while_stage_0_8;
  assign input_mem_banks_read_1_read_data_and_cse = PECoreRun_wen & and_525_cse;
  assign input_mem_banks_read_1_read_data_and_5_enex5 = input_mem_banks_read_1_read_data_and_cse
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  assign weight_mem_run_3_for_5_and_177_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_175_cse = reg_weight_mem_run_3_for_5_and_162_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_176_cse = reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_178_cse = reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_179_cse = reg_weight_mem_run_3_for_5_and_166_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_181_cse = reg_weight_mem_run_3_for_5_and_168_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_188_cse = reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_185_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_189_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign or_691_cse = (~ weight_mem_run_3_for_land_1_lpi_1_dfm_2) | PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  assign or_687_cse = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  assign weight_port_read_out_data_and_enex5 = PECoreRun_wen & (~(or_dcpl_219 | (~
      weight_mem_run_3_for_land_2_lpi_1_dfm_3))) & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000000;
  assign weight_mem_run_3_for_aelse_and_cse = PECoreRun_wen & while_stage_0_7;
  assign weight_port_read_out_data_and_1_cse = PECoreRun_wen & (~(or_dcpl_219 | (~
      weight_mem_run_3_for_land_3_lpi_1_dfm_3)));
  assign weight_port_read_out_data_and_79_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000000;
  assign data_in_tmp_operator_2_for_and_1_cse = PECoreRun_wen & and_dcpl_48 & weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  assign weight_port_read_out_data_and_80_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000001;
  assign weight_port_read_out_data_and_81_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000002;
  assign weight_port_read_out_data_and_82_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000003;
  assign weight_port_read_out_data_and_83_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000004;
  assign weight_port_read_out_data_and_84_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000005;
  assign weight_port_read_out_data_and_85_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000006;
  assign PECore_RunMac_if_and_4_cse = PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & rva_in_reg_rw_sva_st_1_5)) & while_stage_0_7;
  assign rva_in_reg_rw_and_2_cse = PECoreRun_wen & and_dcpl_59;
  assign input_mem_banks_read_1_read_data_and_1_enex5 = PECoreRun_wen & reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  assign PECore_RunMac_if_and_5_cse = PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign nor_419_cse = ~((weight_read_addrs_7_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_288_nl = MUX_s_1_2_2((weight_read_addrs_7_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_7_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_7_lpi_1_dfm_3_2_0[0]);
  assign mux_289_cse = MUX_s_1_2_2(mux_288_nl, nor_419_cse, weight_read_addrs_7_lpi_1_dfm_3_2_0[2]);
  assign and_1053_cse = (mux_289_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign and_1062_cse = (and_1053_cse | or_dcpl_336 | or_dcpl_325) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7 & PECoreRun_wen;
  assign and_1066_cse = (((((weight_read_addrs_7_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[2])) | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2) | or_dcpl_336 | PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7 & PECoreRun_wen;
  assign xor_5_cse = (weight_read_addrs_5_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_5_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign and_1085_cse = (xor_5_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign and_1086_cse = (and_1085_cse | weight_mem_run_3_for_5_and_95_itm_2 | weight_mem_run_3_for_5_and_94_itm_2
      | weight_mem_run_3_for_5_and_92_itm_2) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7 & PECoreRun_wen;
  assign nor_425_cse = ~((weight_read_addrs_5_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_300_nl = MUX_s_1_2_2((weight_read_addrs_5_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_5_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_5_lpi_1_dfm_3_2_0[0]);
  assign mux_301_nl = MUX_s_1_2_2(mux_300_nl, nor_425_cse, weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign and_1090_cse = (((mux_301_nl | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2) | or_dcpl_368 | weight_mem_run_3_for_5_and_92_itm_2
      | weight_mem_run_3_for_5_and_88_itm_1) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7 & PECoreRun_wen;
  assign weight_mem_run_3_for_aelse_and_4_cse = PECoreRun_wen & while_stage_0_6;
  assign weight_port_read_out_data_3_7_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[111:96]), weight_port_read_out_data_3_7_sva_dfm_1,
      {weight_mem_run_3_for_5_and_166 , weight_mem_run_3_for_5_asn_306 , weight_mem_run_3_for_5_asn_308
      , weight_mem_run_3_for_5_and_28_itm_1 , weight_mem_run_3_for_5_asn_310 , reg_weight_mem_run_3_for_5_and_30_itm_2_cse
      , weight_mem_run_3_for_5_and_31_itm_1 , weight_mem_run_3_for_5_asn_312 , (~
      weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign xor_13_cse = (weight_read_addrs_3_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_3_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_3_lpi_1_dfm_3_2_0[2]);
  assign and_1118_cse = (xor_13_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_port_read_out_data_3_6_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[95:80]), weight_port_read_out_data_3_6_sva_dfm_1,
      {weight_mem_run_3_for_5_and_166 , weight_mem_run_3_for_5_asn_306 , weight_mem_run_3_for_5_asn_308
      , reg_weight_mem_run_3_for_5_and_20_itm_2_cse , weight_mem_run_3_for_5_asn_310
      , weight_mem_run_3_for_5_and_22_itm_1 , weight_mem_run_3_for_5_and_31_itm_1
      , weight_mem_run_3_for_5_asn_312 , (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign weight_port_read_out_data_3_5_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[79:64]), weight_port_read_out_data_3_5_sva_dfm_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse , weight_mem_run_3_for_5_asn_306
      , weight_mem_run_3_for_5_asn_308 , reg_weight_mem_run_3_for_5_and_20_itm_2_cse
      , weight_mem_run_3_for_5_asn_310 , reg_weight_mem_run_3_for_5_and_30_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , weight_mem_run_3_for_5_asn_312
      , (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign weight_port_read_out_data_3_4_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[63:48]), weight_port_read_out_data_3_4_sva_dfm_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse , weight_mem_run_3_for_5_asn_306
      , weight_mem_run_3_for_5_asn_308 , reg_weight_mem_run_3_for_5_and_20_itm_2_cse
      , weight_mem_run_3_for_5_asn_310 , reg_weight_mem_run_3_for_5_and_30_itm_2_cse
      , weight_mem_run_3_for_5_and_31_itm_1 , weight_mem_run_3_for_5_and_8_itm_1
      , (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign nor_428_cse = ~((weight_read_addrs_3_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign weight_read_addrs_and_3_cse = PECoreRun_wen & ((weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
      & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]))) | ((~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]))
      & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1))
      & and_dcpl_71;
  assign weight_read_addrs_and_enex5 = weight_read_addrs_and_3_cse & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse = PECoreRun_wen & and_dcpl_80;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse
      & (reg_weight_read_addrs_6_14_1_lpi_1_dfm_1_enexo | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1);
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse = PECoreRun_wen & and_dcpl_82;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse
      & (reg_weight_read_addrs_6_14_1_lpi_1_dfm_1_enexo_1 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo_1
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1
      | reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1);
  assign while_if_and_11_cse = PECoreRun_wen & while_stage_0_5;
  assign weight_mem_read_arbxbar_arbiters_next_and_cse = accum_vector_data_and_cse
      & ((nor_cse & nor_197_cse & nor_198_cse & nor_199_cse) | or_dcpl_60);
  assign weight_mem_read_arbxbar_arbiters_next_and_53_cse = accum_vector_data_and_cse
      & (and_108_cse | or_dcpl_60);
  assign weight_mem_read_arbxbar_arbiters_next_and_59_cse = accum_vector_data_and_cse
      & or_dcpl_63;
  assign weight_mem_read_arbxbar_arbiters_next_and_65_cse = accum_vector_data_and_cse
      & or_dcpl_64;
  assign weight_mem_read_arbxbar_arbiters_next_and_71_cse = accum_vector_data_and_cse
      & or_187_cse;
  assign weight_mem_read_arbxbar_arbiters_next_and_77_cse = accum_vector_data_and_cse
      & (and_129_cse | or_dcpl_60);
  assign weight_mem_read_arbxbar_arbiters_next_and_83_cse = accum_vector_data_and_cse
      & (and_dcpl_136 | or_dcpl_60);
  assign weight_mem_read_arbxbar_arbiters_next_and_89_cse = accum_vector_data_and_cse
      & ((~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4));
  assign weight_read_addrs_and_5_cse = PECoreRun_wen & (and_dcpl_144 | and_dcpl_143
      | and_dcpl_142 | and_dcpl_141 | and_dcpl_140 | and_dcpl_139 | and_dcpl_138
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | and_dcpl_137) & while_stage_0_4;
  assign weight_write_data_data_and_cse = PECoreRun_wen & ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7:6]!=2'b00))
      & and_dcpl_146;
  assign weight_write_data_data_and_24_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_25_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_26_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_27_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_28_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_29_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_30_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_31_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_addrs_and_enex5 = weight_write_data_data_and_cse & reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  assign weight_mem_write_arbxbar_xbar_for_1_for_and_cse = PECoreRun_wen & and_dcpl_146;
  assign mux_29_nl = MUX_s_1_2_2(mux_tmp_16, mux_tmp_13, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1);
  assign mux_30_nl = MUX_s_1_2_2(mux_tmp_27, mux_29_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign while_mux_1276_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_17_nl = MUX_s_1_2_2(mux_tmp_16, mux_tmp_13, while_mux_1276_nl);
  assign mux_28_nl = MUX_s_1_2_2(mux_tmp_27, mux_17_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign mux_31_nl = MUX_s_1_2_2(mux_30_nl, mux_28_nl, while_stage_0_5);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
      = PECoreRun_wen & mux_31_nl & and_dcpl_154;
  assign weight_read_addrs_and_7_cse = PECoreRun_wen & and_dcpl_154;
  assign PECore_RunFSM_switch_lp_and_cse = PECoreRun_wen & while_stage_0_4;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 & and_dcpl_154;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 & and_dcpl_154;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13 & and_dcpl_154;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14 & and_dcpl_154;
  assign Arbiter_8U_Roundrobin_pick_1_and_15_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8
      & and_dcpl_154;
  assign Arbiter_8U_Roundrobin_pick_and_cse = PECoreRun_wen & (while_stage_0_4 |
      and_dcpl_582) & fsm_output & or_dcpl_60;
  assign Arbiter_8U_Roundrobin_pick_1_and_22_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9
      & and_dcpl_154;
  assign Arbiter_8U_Roundrobin_pick_1_and_64_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign weight_write_data_data_and_8_cse = PECoreRun_wen & and_dcpl_189;
  assign weight_write_data_data_and_32_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_33_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_34_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_35_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_36_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_37_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_38_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_39_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  assign weight_write_addrs_and_3_enex5 = weight_write_data_data_and_8_cse & reg_weight_write_addrs_lpi_1_dfm_1_1_enexo;
  assign rva_in_reg_rw_and_3_cse = PECoreRun_wen & while_stage_0_3;
  assign weight_read_addrs_and_29_enex5 = weight_write_data_data_and_8_cse & reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  assign state_and_cse = accum_vector_data_and_cse & nand_58_cse;
  assign nor_431_cse = ~((~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1);
  assign pe_config_num_manager_and_cse = PECoreRun_wen & (~(or_dcpl_233 | or_dcpl_231
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]))));
  assign rva_in_reg_rw_and_4_cse = PECoreRun_wen & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign PECore_UpdateFSM_switch_lp_and_11_cse = PECoreRun_wen & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign or_804_cse = (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_1331_cse = pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
      & PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
  assign pe_config_UpdateManagerCounter_if_if_and_enex5 = PECoreRun_wen & reg_pe_config_num_output_enexo;
  assign nor_438_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:10]!=2'b00));
  assign and_1173_cse = (((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:2]==8'b00000000)
      & nor_438_cse & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:12]!=2'b00)))
      & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:14]!=2'b00))) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | (~(reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3))) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01)
      & rva_in_PopNB_mioi_return_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]==2'b00)
      & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & rva_in_reg_rw_and_4_cse;
  assign PECore_DecodeAxiRead_switch_lp_and_cse = PECoreRun_wen & (~(nand_58_cse
      | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
  assign PECore_DecodeAxiWrite_switch_lp_and_cse = PECoreRun_wen & (~ or_dcpl_231);
  assign and_1178_nl = ((~ while_stage_0_10) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8)
      & or_tmp_374;
  assign and_1177_nl = (PECore_RunMac_PECore_RunMac_if_and_svs_8 | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_8)
      | (~ while_stage_0_10) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8)
      & or_tmp_374;
  assign or_814_nl = (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8) | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
  assign mux_315_nl = MUX_s_1_2_2(and_1178_nl, and_1177_nl, or_814_nl);
  assign and_1179_cse = mux_315_nl & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9)
      & rva_in_reg_rw_and_cse;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_or_1_cse = ((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3==3'b010)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3) | ((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3==3'b100)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_929_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_28 & (~ or_dcpl);
  assign and_930_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_35 & (~ or_dcpl);
  assign and_931_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_1_cse & (~ or_dcpl);
  assign and_932_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1
      & (~ or_dcpl);
  assign and_933_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      & (~ or_dcpl);
  assign and_934_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1
      & (~ or_dcpl);
  assign and_935_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1
      & (~ or_dcpl);
  assign nor_397_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl);
  assign weight_read_addrs_and_16_cse = PECoreRun_wen & weight_mem_run_3_for_land_5_lpi_1_dfm_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign weight_port_read_out_data_and_28_cse = PECoreRun_wen & ((weight_mem_run_3_for_land_1_lpi_1_dfm_3
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5))
      | while_and_30_tmp) & while_stage_0_7;
  assign weight_port_read_out_data_and_32_cse = PECoreRun_wen & (~(or_dcpl_222 |
      (~ weight_mem_run_3_for_land_7_lpi_1_dfm_2)));
  assign weight_port_read_out_data_and_40_cse = PECoreRun_wen & (~(or_dcpl_222 |
      (~ weight_mem_run_3_for_land_2_lpi_1_dfm_2)));
  assign weight_port_read_out_data_and_48_cse = PECoreRun_wen & (~(or_dcpl_222 |
      (~ weight_mem_run_3_for_land_5_lpi_1_dfm_2)));
  assign or_17_nl = (~ weight_mem_run_3_for_weight_mem_run_3_for_and_3_tmp) | (~
      while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign or_16_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_run_3_for_land_4_lpi_1_dfm_1);
  assign mux_3_nl = MUX_s_1_2_2(or_17_nl, or_16_nl, while_stage_0_6);
  assign weight_port_read_out_data_and_68_cse = PECoreRun_wen & (~(or_dcpl_222 |
      (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2) | (~ fsm_output))) & mux_3_nl;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_4_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_103_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_108_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_2_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_109_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse = PECoreRun_wen & weight_mem_run_3_for_land_1_lpi_1_dfm_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign weight_read_addrs_and_19_cse = PECoreRun_wen & and_dcpl_78;
  assign and_739_cse = (reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign or_187_cse = (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp);
  assign and_741_cse = (~((~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp)
      | nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_1_tmp))
      | Arbiter_8U_Roundrobin_pick_1_if_1_and_8_tmp | Arbiter_8U_Roundrobin_pick_1_if_1_and_5_tmp;
  assign and_742_cse = (~ nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_1_tmp)
      & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
  assign and_740_cse = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) & weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp;
  assign mux_256_cse = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp,
      and_733_cse, weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_24_cse
      = accum_vector_data_and_cse & or_dcpl_60;
  assign weight_read_addrs_and_30_enex5 = weight_write_data_data_and_8_cse & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  assign operator_15_false_1_and_cse = PECoreRun_wen & (~(and_dcpl_580 | or_dcpl_60));
  assign PEManager_15U_PEManagerWrite_and_enex5 = PECoreRun_wen & reg_rva_in_reg_rw_sva_st_1_1_cse
      & (~ PECore_DecodeAxiWrite_switch_lp_nor_tmp_1) & PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1
      & (~ PECore_DecodeAxiWrite_switch_lp_equal_tmp_2) & (~ PECore_DecodeAxiWrite_switch_lp_equal_tmp_1)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_in_reg_data_sva_1_enexo;
  assign pe_manager_num_input_and_cse = PECoreRun_wen & (~(or_dcpl_233 | nand_58_cse
      | or_dcpl_273));
  assign pe_config_is_valid_and_cse = PECoreRun_wen & (~(PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1
      | PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (~ nand_58_cse);
  assign while_if_and_15_cse = PECoreRun_wen & and_dcpl_197;
  assign rva_in_reg_rw_and_5_cse = PECoreRun_wen & and_dcpl_71;
  assign rva_in_reg_rw_and_6_cse = PECoreRun_wen & and_dcpl_237;
  assign input_mem_banks_read_read_data_and_9_cse = PECoreRun_wen & and_dcpl_241
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6) & input_read_req_valid_lpi_1_dfm_1_8;
  assign input_mem_banks_read_read_data_and_52_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_53_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_54_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_55_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse = PECoreRun_wen & and_dcpl_237
      & (~(rva_in_reg_rw_sva_st_1_8 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6))
      & (~(rva_in_reg_rw_sva_8 | input_read_req_valid_lpi_1_dfm_1_8)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  assign PECore_UpdateFSM_switch_lp_and_17_cse = PECoreRun_wen & and_dcpl_45;
  assign input_mem_banks_read_1_read_data_and_2_enex5 = PECoreRun_wen & PECore_RunMac_PECore_RunMac_if_and_svs_st_3
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  assign input_read_req_valid_and_1_cse = PECoreRun_wen & and_dcpl_241;
  assign PECore_DecodeAxiRead_switch_lp_and_7_cse = PECoreRun_wen & and_dcpl_252;
  assign rva_out_reg_data_and_30_cse = PECoreRun_wen & and_dcpl_252 & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_8
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8))
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 & (~ rva_in_reg_rw_sva_st_8);
  assign rva_out_reg_data_and_124_enex5 = rva_out_reg_data_and_30_cse & reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_125_enex5 = rva_out_reg_data_and_30_cse & reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_126_enex5 = rva_out_reg_data_and_30_cse & reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  assign weight_port_read_out_data_and_72_cse = PECoreRun_wen & and_dcpl_237 & (~
      rva_in_reg_rw_sva_st_1_8) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  assign weight_port_read_out_data_and_86_enex5 = weight_port_read_out_data_and_72_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo;
  assign rva_out_reg_data_and_127_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_128_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_129_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_130_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_62_48_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_131_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_127_112_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_132_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_111_96_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_133_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_95_80_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_134_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_79_64_sva_dfm_4_3_enexo;
  assign weight_mem_banks_load_store_for_else_and_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1 & and_dcpl_59;
  assign weight_mem_banks_load_store_for_else_and_24_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1 & and_dcpl_59;
  assign or_202_cse = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2:1]!=2'b00);
  assign nor_275_cse = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2:1]!=2'b00));
  assign and_915_cse = (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]) & nor_275_cse;
  assign and_916_cse = (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]) & and_dcpl_643;
  assign or_639_tmp = and_dcpl_724 | and_916_cse | and_915_cse;
  assign weight_mem_banks_load_store_for_else_and_27_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_mem_banks_load_store_for_else_and_28_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign or_641_nl = and_915_cse | and_916_cse | nor_tmp_191;
  assign mux_259_tmp = MUX_s_1_2_2(nor_tmp_191, or_641_nl, and_dcpl_266);
  assign weight_read_addrs_and_24_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse
      & and_dcpl_279;
  assign and_289_cse = PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]);
  assign rva_in_reg_rw_and_9_cse = PECoreRun_wen & and_dcpl_297;
  assign pe_manager_base_weight_and_5_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse
      & and_dcpl_279;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_117_cse = PECoreRun_wen
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | weight_mem_run_3_for_weight_mem_run_3_for_and_3_tmp) & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_122_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_83_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_89_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_1_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign input_mem_banks_read_read_data_and_18_cse = PECoreRun_wen & and_dcpl_325
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5) & input_read_req_valid_lpi_1_dfm_1_7;
  assign input_mem_banks_read_read_data_and_56_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_57_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_58_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_59_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse = PECoreRun_wen & and_dcpl_297
      & (~(rva_in_reg_rw_sva_st_1_7 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5))
      & (~(input_read_req_valid_lpi_1_dfm_1_7 | rva_in_reg_rw_sva_7)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
  assign PECore_UpdateFSM_switch_lp_and_18_cse = PECoreRun_wen & and_dcpl_48;
  assign input_mem_banks_read_1_read_data_and_3_enex5 = PECoreRun_wen & PECore_RunMac_PECore_RunMac_if_and_svs_st_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  assign or_253_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_125_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp;
  assign or_260_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp;
  assign input_read_req_valid_and_2_cse = PECoreRun_wen & and_dcpl_325;
  assign PECore_DecodeAxiRead_switch_lp_and_11_cse = PECoreRun_wen & and_dcpl_354;
  assign rva_out_reg_data_and_43_cse = PECoreRun_wen & and_dcpl_354 & (~ rva_in_reg_rw_sva_st_7)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_7)
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7));
  assign rva_out_reg_data_and_135_enex5 = rva_out_reg_data_and_43_cse & reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_136_enex5 = rva_out_reg_data_and_43_cse & reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_137_enex5 = rva_out_reg_data_and_43_cse & reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  assign weight_port_read_out_data_and_74_cse = PECoreRun_wen & and_dcpl_297 & (~
      rva_in_reg_rw_sva_st_1_7) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  assign weight_port_read_out_data_and_87_enex5 = weight_port_read_out_data_and_74_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  assign rva_out_reg_data_and_138_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_139_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_140_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_141_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_62_48_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_142_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_127_112_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_143_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_111_96_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_144_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_95_80_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_145_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_79_64_sva_dfm_4_2_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp;
  assign weight_mem_write_arbxbar_xbar_for_empty_and_enex5 = rva_in_reg_rw_and_5_cse
      & reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  assign PECore_RunMac_if_and_7_cse = PECoreRun_wen & and_628_cse;
  assign rva_in_reg_rw_and_12_cse = PECoreRun_wen & and_dcpl_362;
  assign input_mem_banks_read_read_data_and_27_cse = PECoreRun_wen & and_dcpl_365
      & input_read_req_valid_lpi_1_dfm_1_6 & and_dcpl_362;
  assign input_mem_banks_read_read_data_and_60_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_61_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_62_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_63_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse = PECoreRun_wen & and_dcpl_365
      & (~(rva_in_reg_rw_sva_6 | input_read_req_valid_lpi_1_dfm_1_6)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5
      & while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  assign and_374_cse = PECore_UpdateFSM_switch_lp_equal_tmp_3_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign input_read_req_valid_and_3_cse = PECoreRun_wen & (~ rva_in_reg_rw_sva_st_1_6)
      & while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  assign PECore_DecodeAxiRead_switch_lp_and_15_cse = PECoreRun_wen & and_dcpl_379
      & (~ input_read_req_valid_lpi_1_dfm_1_6) & while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  assign rva_out_reg_data_and_54_cse = PECoreRun_wen & and_dcpl_379 & (~ input_read_req_valid_lpi_1_dfm_1_6)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6)
      & (~(rva_in_reg_rw_sva_st_6 | PECore_DecodeAxiRead_switch_lp_nor_tmp_6 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6))
      & and_dcpl_362;
  assign rva_out_reg_data_and_146_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_30_25_sva_dfm_4_enexo;
  assign rva_out_reg_data_and_147_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_23_17_sva_dfm_4_enexo;
  assign rva_out_reg_data_and_148_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_15_9_sva_dfm_6_enexo;
  assign weight_port_read_out_data_and_76_cse = PECoreRun_wen & (~ rva_in_reg_rw_sva_st_1_6)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 & and_dcpl_362;
  assign rva_out_reg_data_and_149_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_150_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_151_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_152_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_62_48_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_153_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_127_112_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_154_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_111_96_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_155_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_95_80_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_156_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_79_64_sva_dfm_4_1_enexo;
  assign rva_in_reg_rw_and_15_cse = PECoreRun_wen & and_dcpl_212;
  assign input_mem_banks_read_read_data_and_36_cse = PECoreRun_wen & and_dcpl_393
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1;
  assign input_mem_banks_read_read_data_and_64_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  assign input_mem_banks_read_read_data_and_65_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1;
  assign input_mem_banks_read_read_data_and_66_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2;
  assign input_mem_banks_read_read_data_and_67_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse = PECoreRun_wen & and_dcpl_212
      & (~(rva_in_reg_rw_sva_st_1_5 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3))
      & (~ rva_in_reg_rw_sva_5) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 &
      (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1);
  assign input_read_req_valid_and_4_cse = PECoreRun_wen & and_dcpl_393;
  assign PECore_DecodeAxiRead_switch_lp_and_19_cse = PECoreRun_wen & and_dcpl_393
      & and_dcpl_400 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1);
  assign rva_out_reg_data_and_65_cse = PECoreRun_wen & and_dcpl_393 & and_dcpl_400
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_5) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4
      & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5) & (~ rva_in_reg_rw_sva_st_5)
      & (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5));
  assign rva_out_reg_data_and_157_enex5 = rva_out_reg_data_and_65_cse & reg_rva_out_reg_data_30_25_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_158_enex5 = rva_out_reg_data_and_65_cse & reg_rva_out_reg_data_23_17_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_159_enex5 = rva_out_reg_data_and_65_cse & reg_rva_out_reg_data_15_9_sva_dfm_5_enexo;
  assign and_1235_cse = (~(((~(rva_in_reg_rw_sva_6 | (~ while_stage_0_8) | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)) | rva_in_reg_rw_sva_st_1_5)
      & rva_in_reg_rw_sva_5)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & PECoreRun_wen & while_stage_0_7;
  assign rva_out_reg_data_and_72_cse = PECoreRun_wen & (~ mux_tmp) & while_stage_0_7;
  assign and_1252_cse = (~ rva_in_reg_rw_sva_6) & while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & fsm_output & (rva_in_reg_rw_sva_5 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      | (~ while_stage_0_7)) & PECoreRun_wen;
  assign rva_out_reg_data_and_80_cse = PECoreRun_wen & not_tmp_147 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign rva_out_reg_data_and_160_enex5 = rva_out_reg_data_and_80_cse & reg_rva_out_reg_data_46_40_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_161_enex5 = rva_out_reg_data_and_80_cse & reg_rva_out_reg_data_39_36_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_162_enex5 = rva_out_reg_data_and_80_cse & reg_rva_out_reg_data_35_32_sva_dfm_1_4_enexo;
  assign nand_58_cse = ~(rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse);
  assign or_868_nl = rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | nand_58_cse;
  assign or_867_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign mux_317_nl = MUX_s_1_2_2(or_868_nl, or_867_nl, while_stage_0_3);
  assign or_866_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | reg_rva_in_reg_rw_sva_2_cse;
  assign mux_318_nl = MUX_s_1_2_2(mux_317_nl, or_866_nl, while_stage_0_4);
  assign or_865_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | rva_in_reg_rw_sva_3;
  assign mux_319_nl = MUX_s_1_2_2(mux_318_nl, or_865_nl, while_stage_0_5);
  assign or_864_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | rva_in_reg_rw_sva_4;
  assign mux_320_nl = MUX_s_1_2_2(mux_319_nl, or_864_nl, while_stage_0_6);
  assign and_1272_cse = mux_320_nl & fsm_output & while_stage_0_7 & PECoreRun_wen
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~ rva_in_reg_rw_sva_5);
  assign nor_472_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_21_cse = PECoreRun_wen & (~ or_tmp_54)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign PECore_DecodeAxiRead_switch_lp_and_23_cse = PECoreRun_wen & (~(or_tmp_54
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
      & while_stage_0_6;
  assign rva_out_reg_data_and_87_cse = PECoreRun_wen & not_tmp_147 & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_4)
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)) & (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1
      | rva_in_reg_rw_sva_st_4)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 &
      and_dcpl_59;
  assign rva_out_reg_data_and_163_enex5 = rva_out_reg_data_and_87_cse & reg_rva_out_reg_data_30_25_sva_dfm_2_enexo;
  assign rva_out_reg_data_and_164_enex5 = rva_out_reg_data_and_87_cse & reg_rva_out_reg_data_23_17_sva_dfm_2_enexo;
  assign rva_out_reg_data_and_165_enex5 = rva_out_reg_data_and_87_cse & reg_rva_out_reg_data_15_9_sva_dfm_4_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse = PECoreRun_wen & and_dcpl_438
      & (~(input_read_req_valid_lpi_1_dfm_1_3 | rva_in_reg_rw_sva_3)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse = PECoreRun_wen & and_dcpl_443
      & (~ rva_in_reg_rw_sva_3) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign input_mem_banks_read_read_data_and_46_enex5 = PECoreRun_wen & and_dcpl_438
      & input_read_req_valid_lpi_1_dfm_1_3 & and_dcpl_71 & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo;
  assign nor_251_nl = ~(rva_in_reg_rw_sva_3 | input_read_req_valid_lpi_1_dfm_1_3
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1);
  assign mux_91_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, nor_251_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign PECore_DecodeAxiRead_switch_lp_and_27_cse = PECoreRun_wen & mux_91_nl &
      while_stage_0_5;
  assign rva_out_reg_data_and_90_cse = PECoreRun_wen & and_dcpl_443 & (~(rva_in_reg_rw_sva_3
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_3)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3
      | rva_in_reg_rw_sva_st_3)) & and_dcpl_71;
  assign rva_out_reg_data_and_166_enex5 = rva_out_reg_data_and_90_cse & reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_167_enex5 = rva_out_reg_data_and_90_cse & reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_168_enex5 = rva_out_reg_data_and_90_cse & reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_169_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_170_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_171_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_172_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse
      & reg_rva_out_reg_data_62_48_sva_dfm_1_3_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse = PECoreRun_wen & and_dcpl_461
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 & and_dcpl_146;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse = PECoreRun_wen & and_dcpl_461
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign input_mem_banks_read_read_data_and_47_enex5 = PECoreRun_wen & and_dcpl_468
      & input_read_req_valid_lpi_1_dfm_1_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1;
  assign rva_out_reg_data_and_97_cse = PECoreRun_wen & and_dcpl_468 & (~(input_read_req_valid_lpi_1_dfm_1_2
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_2)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1
      & (~(reg_rva_in_reg_rw_sva_2_cse | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign rva_out_reg_data_and_173_enex5 = rva_out_reg_data_and_97_cse & reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  assign rva_out_reg_data_and_174_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_175_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_176_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_177_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse
      & reg_rva_out_reg_data_62_48_sva_dfm_1_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_35_cse = PECoreRun_wen & mux_tmp_92
      & and_dcpl_482;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_36_cse = PECoreRun_wen & and_dcpl_482;
  assign rva_out_reg_data_and_104_enex5 = PECoreRun_wen & (~(input_read_req_valid_lpi_1_dfm_1_1
      | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[0])))
      & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[3:1]==3'b010)
      & and_dcpl_488 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_178_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_36_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_179_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_36_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_180_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_36_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_181_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_36_cse
      & reg_pe_manager_base_input_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_40_cse = PECoreRun_wen & mux_tmp_92
      & and_dcpl_481 & (~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1) &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse = PECoreRun_wen & and_dcpl_204
      & and_dcpl_208 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_45_cse = PECoreRun_wen & and_dcpl_292
      & (~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])))
      & nand_17_cse;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_49_cse = PECoreRun_wen & (or_dcpl_132
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]!=2'b10)) & and_dcpl_238;
  assign PECore_RunScale_and_14_nl = (~ PECore_RunScale_if_for_1_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign PECore_RunScale_and_15_nl = PECore_RunScale_if_for_1_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign act_port_reg_data_31_0_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_31_0_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_24 , PECore_RunScale_and_14_nl , PECore_RunScale_and_15_nl});
  assign PECore_RunScale_and_12_nl = (~ PECore_RunScale_if_for_2_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign PECore_RunScale_and_13_nl = PECore_RunScale_if_for_2_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign act_port_reg_data_63_32_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_63_32_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_24 , PECore_RunScale_and_12_nl , PECore_RunScale_and_13_nl});
  assign PECore_RunScale_and_10_nl = (~ PECore_RunScale_if_for_3_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign PECore_RunScale_and_11_nl = PECore_RunScale_if_for_3_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign act_port_reg_data_95_64_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_95_64_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_24 , PECore_RunScale_and_10_nl , PECore_RunScale_and_11_nl});
  assign PECore_RunScale_and_8_nl = (~ PECore_RunScale_if_for_4_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign PECore_RunScale_and_9_nl = PECore_RunScale_if_for_4_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign act_port_reg_data_127_96_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_127_96_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_24 , PECore_RunScale_and_8_nl , PECore_RunScale_and_9_nl});
  assign PECore_RunScale_and_6_nl = (~ PECore_RunScale_if_for_5_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign PECore_RunScale_and_7_nl = PECore_RunScale_if_for_5_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign act_port_reg_data_159_128_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_159_128_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_24 , PECore_RunScale_and_6_nl , PECore_RunScale_and_7_nl});
  assign PECore_RunScale_and_2_nl = (~ PECore_RunScale_if_for_7_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign PECore_RunScale_and_3_nl = PECore_RunScale_if_for_7_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_10);
  assign act_port_reg_data_223_192_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_223_192_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_24 , PECore_RunScale_and_2_nl , PECore_RunScale_and_3_nl});
  assign and_562_cse = while_stage_0_12 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
      & (~ rva_in_reg_rw_sva_st_1_10);
  assign and_567_cse = while_stage_0_12 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10)
      & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10;
  assign weight_port_read_out_data_5_6_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[95:80]), weight_port_read_out_data_5_6_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_298 , weight_mem_run_3_for_5_asn_300
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_302 , weight_mem_run_3_for_5_and_86_itm_1
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_and_88_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_7_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[111:96]), weight_port_read_out_data_5_7_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_298 , weight_mem_run_3_for_5_asn_300
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_302 , weight_mem_run_3_for_5_and_94_itm_2
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_asn_304 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_4_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[63:48]), weight_port_read_out_data_5_4_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_298 , weight_mem_run_3_for_5_asn_300
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_302 , weight_mem_run_3_for_5_and_86_itm_1
      , weight_mem_run_3_for_5_and_71_itm_1 , weight_mem_run_3_for_5_asn_304 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_5_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[79:64]), weight_port_read_out_data_5_5_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_298 , weight_mem_run_3_for_5_asn_300
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_302 , weight_mem_run_3_for_5_and_86_itm_1
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_and_88_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_2_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[31:16]), weight_port_read_out_data_5_2_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_298 , weight_mem_run_3_for_5_asn_300
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_302 , weight_mem_run_3_for_5_and_94_itm_2
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_asn_304 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_3_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[47:32]), weight_port_read_out_data_5_3_sva_dfm_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_298 , weight_mem_run_3_for_5_asn_300
      , weight_mem_run_3_for_5_and_60_itm_1 , weight_mem_run_3_for_5_asn_302 , weight_mem_run_3_for_5_and_86_itm_1
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_asn_304 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_mem_run_3_for_5_and_36_nl = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b011)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_port_read_out_data_5_0_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]),
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9, weight_port_read_out_data_5_0_sva_dfm_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_298 , weight_mem_run_3_for_5_asn_300
      , weight_mem_run_3_for_5_and_36_nl , weight_mem_run_3_for_5_asn_302 , weight_mem_run_3_for_5_and_86_itm_1
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_asn_304 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_1_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[15:0]), weight_port_read_out_data_5_1_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_298 , weight_mem_run_3_for_5_asn_300
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_302 , weight_mem_run_3_for_5_and_86_itm_1
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_and_88_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_mem_run_3_for_5_and_145_nl = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_port_read_out_data_7_6_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[95:80]), weight_port_read_out_data_7_6_sva_dfm_1,
      {weight_mem_run_3_for_5_and_145_nl , weight_mem_run_3_for_5_asn_290 , weight_mem_run_3_for_5_asn_292
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_294 , weight_mem_run_3_for_5_and_150_itm_2
      , PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_7_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[111:96]), weight_port_read_out_data_7_7_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_290 , weight_mem_run_3_for_5_asn_292
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_294 , PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5
      , weight_mem_run_3_for_5_and_159_itm_2 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_4_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[63:48]), weight_port_read_out_data_7_4_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_290 , weight_mem_run_3_for_5_asn_292
      , PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 , weight_mem_run_3_for_5_asn_294
      , weight_mem_run_3_for_5_and_150_itm_2 , weight_mem_run_3_for_5_and_159_itm_2
      , weight_mem_run_3_for_5_asn_296 , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_5_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[79:64]), weight_port_read_out_data_7_5_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_290 , weight_mem_run_3_for_5_asn_292
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_294 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_159_itm_2 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_2_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[31:16]), weight_port_read_out_data_7_2_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_290 , weight_mem_run_3_for_5_asn_292
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_294 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_159_itm_2 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_3_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[47:32]), weight_port_read_out_data_7_3_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_290 , weight_mem_run_3_for_5_asn_292
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_294 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_159_itm_2 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_0_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]),
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9, weight_port_read_out_data_7_0_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_290 , weight_mem_run_3_for_5_asn_292
      , PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 , weight_mem_run_3_for_5_asn_294
      , weight_mem_run_3_for_5_and_150_itm_2 , weight_mem_run_3_for_5_and_159_itm_2
      , weight_mem_run_3_for_5_asn_296 , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_1_sva_dfm_2 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[15:0]), weight_port_read_out_data_7_1_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_290 , weight_mem_run_3_for_5_asn_292
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_294 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_159_itm_2 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign PECore_RunScale_and_nl = (~ PECore_RunScale_if_for_8_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_9 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_9);
  assign PECore_RunScale_and_1_nl = PECore_RunScale_if_for_8_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_9 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_9);
  assign act_port_reg_data_255_224_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_255_224_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_or_cse , PECore_RunScale_and_nl , PECore_RunScale_and_1_nl});
  assign PECore_RunScale_and_4_nl = (~ PECore_RunScale_if_for_6_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_9 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_9);
  assign PECore_RunScale_and_5_nl = PECore_RunScale_if_for_6_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_9 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_9);
  assign act_port_reg_data_191_160_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_191_160_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_or_cse , PECore_RunScale_and_4_nl , PECore_RunScale_and_5_nl});
  assign and_947_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_35 & (~ or_dcpl_316);
  assign and_948_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_1_cse & (~ or_dcpl_316);
  assign and_949_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1
      & (~ or_dcpl_316);
  assign and_950_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1
      & (~ or_dcpl_316);
  assign and_951_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1
      & (~ or_dcpl_316);
  assign and_952_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1
      & (~ or_dcpl_316);
  assign nor_399_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl_316);
  assign PECore_PushAxiRsp_if_else_mux_18_mx0w2 = MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1_1
      = ~((weight_read_addrs_3_lpi_1_dfm_2_2_0!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_mx0w0 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_mx0w0 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign Arbiter_8U_Roundrobin_pick_nand_22_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_21_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1
      & and_dcpl_78;
  assign weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_22_cse , Arbiter_8U_Roundrobin_pick_and_21_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_22_cse , Arbiter_8U_Roundrobin_pick_and_21_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_22_cse , Arbiter_8U_Roundrobin_pick_and_21_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_22_cse , Arbiter_8U_Roundrobin_pick_and_21_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_22_cse , Arbiter_8U_Roundrobin_pick_and_21_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_22_cse , Arbiter_8U_Roundrobin_pick_and_21_cse});
  assign weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign Arbiter_8U_Roundrobin_pick_nand_10_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_15_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1
      & and_dcpl_78;
  assign weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_15_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_15_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_15_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_15_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_15_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_15_cse});
  assign weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_nand_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_23_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_68_nl = weight_mem_read_arbxbar_arbiters_next_5_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_68_nl,
      weight_mem_read_arbxbar_arbiters_next_5_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_69_nl = weight_mem_read_arbxbar_arbiters_next_5_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_69_nl,
      weight_mem_read_arbxbar_arbiters_next_5_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl = weight_mem_read_arbxbar_arbiters_next_5_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl,
      weight_mem_read_arbxbar_arbiters_next_5_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl = weight_mem_read_arbxbar_arbiters_next_5_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl,
      weight_mem_read_arbxbar_arbiters_next_5_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_cse = weight_mem_read_arbxbar_arbiters_next_5_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_cse,
      weight_mem_read_arbxbar_arbiters_next_5_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_73_nl = weight_mem_read_arbxbar_arbiters_next_5_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_73_nl,
      weight_mem_read_arbxbar_arbiters_next_5_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_23_cse});
  assign weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_nand_35_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_35_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_74_nl = weight_mem_read_arbxbar_arbiters_next_4_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_74_nl,
      weight_mem_read_arbxbar_arbiters_next_4_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_35_cse , Arbiter_8U_Roundrobin_pick_and_35_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_nl = weight_mem_read_arbxbar_arbiters_next_4_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_nl,
      weight_mem_read_arbxbar_arbiters_next_4_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_35_cse , Arbiter_8U_Roundrobin_pick_and_35_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_76_nl = weight_mem_read_arbxbar_arbiters_next_4_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_76_nl,
      weight_mem_read_arbxbar_arbiters_next_4_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_35_cse , Arbiter_8U_Roundrobin_pick_and_35_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_77_nl = weight_mem_read_arbxbar_arbiters_next_4_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_77_nl,
      weight_mem_read_arbxbar_arbiters_next_4_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_35_cse , Arbiter_8U_Roundrobin_pick_and_35_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_cse = weight_mem_read_arbxbar_arbiters_next_4_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_cse,
      weight_mem_read_arbxbar_arbiters_next_4_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_35_cse , Arbiter_8U_Roundrobin_pick_and_35_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_79_nl = weight_mem_read_arbxbar_arbiters_next_4_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_79_nl,
      weight_mem_read_arbxbar_arbiters_next_4_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_35_cse , Arbiter_8U_Roundrobin_pick_and_35_cse});
  assign weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_nand_46_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_43_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_80_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_80_nl,
      weight_mem_read_arbxbar_arbiters_next_3_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_46_cse , Arbiter_8U_Roundrobin_pick_and_43_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_81_nl = weight_mem_read_arbxbar_arbiters_next_3_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_81_nl,
      weight_mem_read_arbxbar_arbiters_next_3_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_46_cse , Arbiter_8U_Roundrobin_pick_and_43_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_82_nl = weight_mem_read_arbxbar_arbiters_next_3_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_82_nl,
      weight_mem_read_arbxbar_arbiters_next_3_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_46_cse , Arbiter_8U_Roundrobin_pick_and_43_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_83_nl = weight_mem_read_arbxbar_arbiters_next_3_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_83_nl,
      weight_mem_read_arbxbar_arbiters_next_3_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_46_cse , Arbiter_8U_Roundrobin_pick_and_43_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_84_nl = weight_mem_read_arbxbar_arbiters_next_3_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_84_nl,
      weight_mem_read_arbxbar_arbiters_next_3_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_46_cse , Arbiter_8U_Roundrobin_pick_and_43_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_85_nl = weight_mem_read_arbxbar_arbiters_next_3_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_85_nl,
      weight_mem_read_arbxbar_arbiters_next_3_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_46_cse , Arbiter_8U_Roundrobin_pick_and_43_cse});
  assign weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_nand_58_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_49_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl = weight_mem_read_arbxbar_arbiters_next_2_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl,
      weight_mem_read_arbxbar_arbiters_next_2_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_58_cse , Arbiter_8U_Roundrobin_pick_and_49_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl = weight_mem_read_arbxbar_arbiters_next_2_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl,
      weight_mem_read_arbxbar_arbiters_next_2_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_58_cse , Arbiter_8U_Roundrobin_pick_and_49_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl = weight_mem_read_arbxbar_arbiters_next_2_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl,
      weight_mem_read_arbxbar_arbiters_next_2_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_58_cse , Arbiter_8U_Roundrobin_pick_and_49_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl = weight_mem_read_arbxbar_arbiters_next_2_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl,
      weight_mem_read_arbxbar_arbiters_next_2_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_58_cse , Arbiter_8U_Roundrobin_pick_and_49_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl,
      weight_mem_read_arbxbar_arbiters_next_2_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_58_cse , Arbiter_8U_Roundrobin_pick_and_49_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl = weight_mem_read_arbxbar_arbiters_next_2_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl,
      weight_mem_read_arbxbar_arbiters_next_2_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_58_cse , Arbiter_8U_Roundrobin_pick_and_49_cse});
  assign weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_nand_70_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_55_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_92_nl = weight_mem_read_arbxbar_arbiters_next_1_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_92_nl,
      weight_mem_read_arbxbar_arbiters_next_1_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_70_cse , Arbiter_8U_Roundrobin_pick_and_55_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl = weight_mem_read_arbxbar_arbiters_next_1_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl,
      weight_mem_read_arbxbar_arbiters_next_1_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_70_cse , Arbiter_8U_Roundrobin_pick_and_55_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl = weight_mem_read_arbxbar_arbiters_next_1_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl,
      weight_mem_read_arbxbar_arbiters_next_1_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_70_cse , Arbiter_8U_Roundrobin_pick_and_55_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_95_nl = weight_mem_read_arbxbar_arbiters_next_1_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_95_nl,
      weight_mem_read_arbxbar_arbiters_next_1_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_70_cse , Arbiter_8U_Roundrobin_pick_and_55_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl,
      weight_mem_read_arbxbar_arbiters_next_1_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_70_cse , Arbiter_8U_Roundrobin_pick_and_55_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_cse = weight_mem_read_arbxbar_arbiters_next_1_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_cse,
      weight_mem_read_arbxbar_arbiters_next_1_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_70_cse , Arbiter_8U_Roundrobin_pick_and_55_cse});
  assign weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_nand_82_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_61_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_98_nl = weight_mem_read_arbxbar_arbiters_next_0_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_98_nl,
      weight_mem_read_arbxbar_arbiters_next_0_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_82_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_99_nl = weight_mem_read_arbxbar_arbiters_next_0_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_99_nl,
      weight_mem_read_arbxbar_arbiters_next_0_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_82_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl = weight_mem_read_arbxbar_arbiters_next_0_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl,
      weight_mem_read_arbxbar_arbiters_next_0_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_82_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl = weight_mem_read_arbxbar_arbiters_next_0_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl,
      weight_mem_read_arbxbar_arbiters_next_0_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_82_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl = weight_mem_read_arbxbar_arbiters_next_0_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl,
      weight_mem_read_arbxbar_arbiters_next_0_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_82_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_103_nl = weight_mem_read_arbxbar_arbiters_next_0_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_103_nl,
      weight_mem_read_arbxbar_arbiters_next_0_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1,
      {and_dcpl_71 , Arbiter_8U_Roundrobin_pick_nand_82_cse , Arbiter_8U_Roundrobin_pick_and_61_cse});
  assign weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_78);
  assign pe_manager_base_weight_sva_mx1_3_0 = MUX_v_4_2_2((pe_manager_base_weight_sva[3:0]),
      (pe_manager_base_weight_sva_dfm_3_1[3:0]), while_stage_0_5);
  assign pe_manager_base_weight_sva_mx2 = MUX_v_15_2_2(pe_manager_base_weight_sva,
      pe_manager_base_weight_sva_dfm_3_1, while_stage_0_5);
  assign nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000001;
  assign PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_1_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000001;
  assign operator_15_false_acc_nl = nl_operator_15_false_acc_nl[13:0];
  assign weight_read_addrs_2_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000011;
  assign PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_3_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_1_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:2])}) + 13'b0000000000001;
  assign operator_15_false_acc_1_nl = nl_operator_15_false_acc_1_nl[12:0];
  assign weight_read_addrs_4_14_2_lpi_1_dfm_1_1 = MUX_v_13_2_2(13'b0000000000000,
      operator_15_false_acc_1_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000101;
  assign PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_5_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_2_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000011;
  assign operator_15_false_acc_2_nl = nl_operator_15_false_acc_2_nl[13:0];
  assign weight_read_addrs_6_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_2_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000111;
  assign PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_7_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112, and_dcpl_580);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97, and_108_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82, and_115_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67, and_122_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign and_645_nl = and_dcpl_636 & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3])));
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52, and_645_nl);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl
      & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37, and_129_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22, and_dcpl_618);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign and_638_nl = (~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])))
      & and_dcpl_625;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7, and_638_nl);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl
      & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1 = (state_2_1_sva[0]) & (~((state_2_1_sva[1])
      | state_0_sva));
  assign state_mux_1_cse = MUX_v_2_2_2(state_2_1_sva, state_2_1_sva_dfm_1, while_stage_0_3);
  assign state_0_sva_mx1 = MUX_s_1_2_2(PECore_UpdateFSM_next_state_0_lpi_1_dfm_4,
      state_0_sva, or_dcpl_226);
  assign while_or_262_nl = (~(PECore_UpdateFSM_switch_lp_equal_tmp_5_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1148_cse_1;
  assign while_and_2_nl = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign pe_config_manager_counter_sva_mx0w0 = MUX1HOT_v_4_3_2(pe_config_manager_counter_sva,
      pe_config_manager_counter_sva_dfm_3_1, pe_config_manager_counter_sva_dfm_1,
      {while_or_262_nl , while_and_2_nl , while_asn_631});
  assign pe_config_manager_counter_sva_mx1 = MUX_v_4_2_2(pe_config_manager_counter_sva,
      pe_config_manager_counter_sva_mx0w0, while_stage_0_3);
  assign PECore_PushOutput_PECore_PushOutput_if_and_svs_1 = (state_mux_1_cse[1])
      & (~((state_mux_1_cse[0]) | state_0_sva_mx1));
  assign PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1 = ~(PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_tmp_129);
  assign pe_config_input_counter_and_cse = while_asn_631 & while_stage_0_3;
  assign nl_operator_8_false_acc_nl = pe_config_input_counter_sva + 8'b00000001;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[7:0];
  assign pe_config_UpdateInputCounter_not_nl = ~ pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl = MUX_v_8_2_2(8'b00000000,
      operator_8_false_acc_nl, pe_config_UpdateInputCounter_not_nl);
  assign pe_config_input_counter_nand_nl = ~(while_stage_0_3 & (~((~(PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1148_cse_1)));
  assign pe_config_input_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_input_counter_sva,
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl, pe_config_input_counter_sva_dfm_1,
      {pe_config_input_counter_nand_nl , and_374_cse , pe_config_input_counter_and_cse});
  assign nl_operator_8_false_1_acc_nl = pe_config_output_counter_sva + 8'b00000001;
  assign operator_8_false_1_acc_nl = nl_operator_8_false_1_acc_nl[7:0];
  assign pe_config_UpdateManagerCounter_if_not_9_nl = ~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl
      = MUX_v_8_2_2(8'b00000000, operator_8_false_1_acc_nl, pe_config_UpdateManagerCounter_if_not_9_nl);
  assign pe_config_output_counter_nand_nl = ~(while_stage_0_3 & (~((~(and_1331_cse
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1148_cse_1)));
  assign while_and_75_nl = and_1331_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign pe_config_output_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_output_counter_sva,
      pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl,
      pe_config_output_counter_sva_dfm_1, {pe_config_output_counter_nand_nl , while_and_75_nl
      , pe_config_input_counter_and_cse});
  assign and_628_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_if_and_2_m1c = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & and_628_cse;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl
      = pe_config_is_zero_first_sva & (~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1);
  assign while_if_or_nl = (~((~((~ PECore_UpdateFSM_switch_lp_equal_tmp_5_1) & and_628_cse))
      & while_stage_0_3)) | ((~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1)
      & while_if_and_2_m1c);
  assign while_if_and_4_nl = pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
      & while_if_and_2_m1c;
  assign pe_config_is_zero_first_sva_mx1 = MUX1HOT_s_1_3_2(while_if_mux_19_itm_1,
      pe_config_is_zero_first_sva, pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl,
      {and_dcpl_189 , while_if_or_nl , while_if_and_4_nl});
  assign PECore_UpdateFSM_switch_lp_equal_tmp_6 = state_0_sva_mx1 & (state_mux_1_cse==2'b00);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1 = (state_mux_1_cse[0])
      & (~((state_mux_1_cse[1]) | state_0_sva_mx1));
  assign pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1
      = ~((pe_config_manager_counter_sva_mx1 != (operator_4_false_acc_sdt_sva_1[3:0]))
      | (operator_4_false_acc_sdt_sva_1[4]));
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18:17]==2'b11)
      & nor_472_cse;
  assign weight_mem_run_3_for_land_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1);
  assign weight_mem_run_3_for_land_6_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1);
  assign weight_mem_run_3_for_weight_mem_run_3_for_and_3_tmp = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2_1);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6,
      or_dcpl_225);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0,
      or_dcpl_225);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5,
      or_dcpl_225);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1,
      or_dcpl_225);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4,
      or_dcpl_225);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2,
      or_dcpl_225);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3,
      or_dcpl_225);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0101);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_3_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_3_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_3_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_125_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  assign weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1_1 = (pe_manager_base_weight_sva[2:0]==3'b111)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1_1 = (pe_manager_base_weight_sva[2:0]==3'b101)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b100)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b010)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b001)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign weight_mem_run_3_for_land_1_lpi_1_dfm_1_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1 = MUX_v_3_2_2(3'b000,
      (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0]), weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp = MUX_s_1_8_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp
      | (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp));
  assign while_and_114_rgt = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_118_rgt = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_122_rgt = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_126_rgt = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_130_rgt = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_134_rgt = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_138_rgt = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_142_rgt = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_146_rgt = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_150_rgt = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_154_rgt = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_158_rgt = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_162_rgt = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_166_rgt = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_170_rgt = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_174_rgt = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_178_rgt = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_182_rgt = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_186_rgt = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_190_rgt = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_194_rgt = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_198_rgt = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_202_rgt = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_206_rgt = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_210_rgt = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_214_rgt = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_218_rgt = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_222_rgt = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_226_rgt = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_230_rgt = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_234_rgt = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_238_rgt = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_242_rgt = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_246_rgt = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_250_rgt = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_254_rgt = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_258_rgt = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_262_rgt = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_266_rgt = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_270_rgt = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_274_rgt = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_278_rgt = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_282_rgt = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_286_rgt = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_290_rgt = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_294_rgt = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_298_rgt = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_302_rgt = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_306_rgt = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_310_rgt = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_314_rgt = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_318_rgt = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_322_rgt = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_326_rgt = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_330_rgt = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_334_rgt = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_338_rgt = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_342_rgt = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_346_rgt = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_350_rgt = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_354_rgt = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_358_rgt = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_362_rgt = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_366_rgt = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_370_rgt = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_374_rgt = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_378_rgt = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_382_rgt = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_386_rgt = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_390_rgt = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_394_rgt = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_398_rgt = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_402_rgt = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_406_rgt = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_410_rgt = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_414_rgt = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_418_rgt = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_422_rgt = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_426_rgt = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_430_rgt = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_434_rgt = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_438_rgt = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_442_rgt = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_446_rgt = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_450_rgt = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_454_rgt = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_458_rgt = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_462_rgt = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_466_rgt = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_470_rgt = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_474_rgt = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_478_rgt = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_482_rgt = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_486_rgt = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_490_rgt = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_494_rgt = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_498_rgt = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_502_rgt = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_506_rgt = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_510_rgt = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_514_rgt = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_518_rgt = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_522_rgt = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_526_rgt = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_530_rgt = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_534_rgt = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_538_rgt = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_542_rgt = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_546_rgt = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_550_rgt = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_554_rgt = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_558_rgt = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_562_rgt = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_566_rgt = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_570_rgt = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_574_rgt = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_578_rgt = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_582_rgt = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_586_rgt = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_590_rgt = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_594_rgt = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_598_rgt = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_602_rgt = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_606_rgt = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_610_rgt = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_614_rgt = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_618_rgt = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_622_rgt = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_626_rgt = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_630_rgt = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_634_rgt = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_638_rgt = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_642_rgt = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_646_rgt = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_650_rgt = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_654_rgt = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_658_rgt = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_662_rgt = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_666_rgt = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_670_rgt = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_674_rgt = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_678_rgt = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_682_rgt = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_686_rgt = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_690_rgt = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_694_rgt = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_698_rgt = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_702_rgt = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_706_rgt = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_710_rgt = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_714_rgt = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_718_rgt = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_722_rgt = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_726_rgt = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_730_rgt = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_734_rgt = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_738_rgt = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_742_rgt = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_746_rgt = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_750_rgt = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_754_rgt = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_758_rgt = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_762_rgt = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_766_rgt = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_770_rgt = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_774_rgt = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_778_rgt = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_782_rgt = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_786_rgt = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_790_rgt = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_794_rgt = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_798_rgt = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_802_rgt = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_806_rgt = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_810_rgt = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_814_rgt = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_818_rgt = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_822_rgt = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_826_rgt = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_830_rgt = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_834_rgt = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_838_rgt = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_842_rgt = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_846_rgt = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_850_rgt = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_854_rgt = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_858_rgt = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_862_rgt = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_866_rgt = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_870_rgt = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_874_rgt = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_878_rgt = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_882_rgt = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_886_rgt = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_890_rgt = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_894_rgt = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_898_rgt = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_902_rgt = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_906_rgt = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_910_rgt = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_914_rgt = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_918_rgt = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_922_rgt = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_926_rgt = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_930_rgt = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_934_rgt = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_938_rgt = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_942_rgt = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_946_rgt = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_950_rgt = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_954_rgt = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_958_rgt = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_962_rgt = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_966_rgt = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_970_rgt = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_974_rgt = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_978_rgt = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_982_rgt = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_986_rgt = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_990_rgt = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_994_rgt = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_998_rgt = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1002_rgt = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1006_rgt = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1010_rgt = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1014_rgt = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1018_rgt = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1022_rgt = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1026_rgt = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1030_rgt = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1034_rgt = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1038_rgt = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1042_rgt = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1046_rgt = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1050_rgt = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1054_rgt = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1058_rgt = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1062_rgt = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1066_rgt = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1070_rgt = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1074_rgt = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1078_rgt = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1082_rgt = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1086_rgt = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1090_rgt = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1094_rgt = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1098_rgt = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1102_rgt = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1106_rgt = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1110_rgt = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1114_rgt = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1118_rgt = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1122_rgt = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1126_rgt = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1130_rgt = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1134_rgt = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign PECore_PushAxiRsp_mux_24_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_5,
      PECore_PushAxiRsp_mux_10_itm_1, rva_in_reg_rw_sva_5);
  assign PECore_PushAxiRsp_if_else_mux_10_mx0w2 = MUX_s_1_2_2(PECore_PushAxiRsp_mux_24_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1);
  assign while_if_while_if_and_16_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_127_112_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_127_112_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_16_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_111_96_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_67
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_17_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_111_96_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_111_96_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_17_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_95_80_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_67
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_18_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_95_80_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_95_80_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_18_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_79_64_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_67
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_19_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_79_64_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_79_64_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_19_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_63_48_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_67
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_62_48_sva_dfm_6_mx1 = MUX_v_15_2_2(rva_out_reg_data_62_48_sva_dfm_4_1,
      rva_out_reg_data_62_48_sva_dfm_6, or_dcpl_279);
  assign rva_out_reg_data_46_40_sva_dfm_6_mx1 = MUX_v_7_2_2(rva_out_reg_data_46_40_sva_dfm_4_1,
      rva_out_reg_data_46_40_sva_dfm_6, or_dcpl_279);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1 = MUX_v_4_2_2(rva_out_reg_data_39_36_sva_dfm_4_1,
      rva_out_reg_data_39_36_sva_dfm_6, or_dcpl_279);
  assign rva_out_reg_data_35_32_sva_dfm_6_mx1 = MUX_v_4_2_2(rva_out_reg_data_35_32_sva_dfm_4_1,
      rva_out_reg_data_35_32_sva_dfm_6, or_dcpl_279);
  assign pe_manager_base_input_sva_mx1 = MUX_v_15_2_2(pe_manager_base_input_sva,
      pe_manager_base_input_sva_dfm_3_1, while_stage_0_3);
  assign PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
      & PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3
      | and_289_cse);
  assign PECore_DecodeAxiRead_switch_lp_nor_tmp_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_RunScale_PECore_RunScale_if_and_1_svs_1 = (state_mux_1_cse[0]) &
      state_0_sva_mx1 & (~ (state_mux_1_cse[1]));
  assign PECore_DecodeAxiRead_switch_lp_nor_9_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 | PECore_DecodeAxiRead_switch_lp_nor_tmp_10);
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1 = ~(input_read_req_valid_lpi_1_dfm_1_10
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign PECore_RunScale_if_for_7_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_5_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_4_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_3_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_2_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_1_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0 = MUX_v_128_2_2(weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0 = MUX_v_112_2_2(weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_16,
      (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:16]), weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_load_store_1_for_else_else_and_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_or_nl = (weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1);
  assign weight_mem_banks_load_store_1_for_else_else_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9 = MUX1HOT_v_16_6_2(BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1,
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1,
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[15:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[15:0]),
      {weight_mem_banks_load_store_1_for_else_else_and_nl , weight_mem_banks_load_store_1_for_else_else_or_nl
      , weight_mem_banks_load_store_1_for_else_else_and_4_nl , weight_mem_banks_load_store_1_for_else_else_and_6_nl
      , weight_mem_banks_load_store_1_for_else_else_and_8_nl , weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2});
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1 = (~(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_sva_1 | mux_144_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_sva_1 & (~ mux_144_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_2_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_sva_1) & not_tmp_388;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_sva_1 & not_tmp_388;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_sva_1) & and_dcpl_674;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_sva_1 & and_dcpl_674;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]),
      {mux_tmp_137 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_2_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_sva_1,
      {mux_tmp_137 , (~ mux_144_itm) , not_tmp_388 , and_dcpl_674});
  assign and_882_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  assign and_881_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  assign and_880_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  assign and_886_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) & while_mux_1329_tmp;
  assign and_885_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) & while_mux_1331_tmp;
  assign and_884_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) & while_mux_1330_tmp;
  assign and_883_cse = weight_mem_read_arbxbar_arbiters_next_7_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign and_887_cse = while_mux_1328_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign nor_384_nl = ~(and_880_cse | and_881_cse | and_882_cse | and_883_cse | or_tmp_141);
  assign nor_385_nl = ~(and_884_cse | and_885_cse | and_886_cse | and_887_cse | or_tmp_139);
  assign mux_159_nl = MUX_s_1_2_2(nor_384_nl, nor_385_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl,
      mux_159_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_6_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1) & not_tmp_393;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 & not_tmp_393;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 | mux_181_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 & (~ mux_181_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1) & and_dcpl_677;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 & and_dcpl_677;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]),
      {mux_tmp_160 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_6_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1,
      {mux_tmp_160 , not_tmp_393 , (~ mux_181_itm) , and_dcpl_677});
  assign and_888_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  assign and_893_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) & while_mux_1319_tmp;
  assign and_891_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  assign and_890_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  assign and_889_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  assign and_896_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & while_mux_1323_tmp;
  assign and_895_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) & while_mux_1321_tmp;
  assign and_894_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & while_mux_1322_tmp;
  assign and_897_cse = while_mux_1324_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign and_892_cse = weight_mem_read_arbxbar_arbiters_next_6_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign nor_386_nl = ~(and_888_cse | and_889_cse | and_890_cse | and_891_cse | and_892_cse
      | or_tmp_177);
  assign nor_387_nl = ~(and_893_cse | and_894_cse | and_895_cse | and_896_cse | and_897_cse
      | or_tmp_175);
  assign mux_189_nl = MUX_s_1_2_2(nor_386_nl, nor_387_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl,
      mux_189_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1) & and_dcpl_680;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 & and_dcpl_680;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1) & and_dcpl_681;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 & and_dcpl_681;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1) & and_dcpl_684;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 & and_dcpl_684;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]),
      {and_dcpl_678 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1,
      {and_dcpl_678 , and_dcpl_680 , and_dcpl_681 , and_dcpl_684});
  assign operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1) & and_dcpl_689;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 & and_dcpl_689;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1) & and_dcpl_690;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 & and_dcpl_690;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1) & and_dcpl_693;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 & and_dcpl_693;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]),
      {and_dcpl_686 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1,
      operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1, {and_dcpl_686 , and_dcpl_689
      , and_dcpl_690 , and_dcpl_693});
  assign operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_24_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1) & and_dcpl_696;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 & and_dcpl_696;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1) & and_dcpl_697;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 & and_dcpl_697;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1) & and_dcpl_703;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 & and_dcpl_703;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]),
      {weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_24_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1,
      operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1, {weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse
      , and_dcpl_696 , and_dcpl_697 , and_dcpl_703});
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse
      = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign and_711_nl = (~ mux_tmp_199) & and_dcpl_695;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse,
      weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl,
      and_711_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 | mux_228_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 & (~ mux_228_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 | mux_241_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 & (~ mux_241_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1) & and_dcpl_705;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 & and_dcpl_705;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]),
      {mux_tmp_215 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1,
      {mux_tmp_215 , (~ mux_228_itm) , (~ mux_241_itm) , and_dcpl_705});
  assign and_903_cse = weight_mem_read_arbxbar_arbiters_next_1_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign and_910_cse = Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign and_904_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  assign and_899_cse = weight_mem_read_arbxbar_arbiters_next_1_5_sva & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign and_901_cse = weight_mem_read_arbxbar_arbiters_next_1_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign and_900_cse = weight_mem_read_arbxbar_arbiters_next_1_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign and_898_cse = weight_mem_read_arbxbar_arbiters_next_1_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign and_906_cse = Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign and_908_cse = Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign and_907_cse = Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign and_905_cse = Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign and_902_cse = weight_mem_read_arbxbar_arbiters_next_1_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign and_909_cse = Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  assign or_613_nl = and_898_cse | and_899_cse | and_900_cse | and_901_cse | and_902_cse
      | and_903_cse | and_904_cse;
  assign or_607_nl = and_905_cse | and_906_cse | and_907_cse | and_908_cse | and_909_cse
      | and_910_cse | nor_tmp_127;
  assign mux_252_nl = MUX_s_1_2_2(or_tmp_304, or_607_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_595_nl = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])
      | nor_tmp_127;
  assign mux_251_nl = MUX_s_1_2_2(or_tmp_304, or_595_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign mux_253_nl = MUX_s_1_2_2(mux_252_nl, mux_251_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_254_nl = MUX_s_1_2_2(or_613_nl, mux_253_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl,
      mux_254_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_mx0w0
      = weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1);
  assign nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_3_mux_mx0w1
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1, weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1) & and_dcpl_711;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 & and_dcpl_711;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1) & and_dcpl_714;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 & and_dcpl_714;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_6_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_mx0w0,
      nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_3_mux_mx0w1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]),
      {and_dcpl_707 , and_dcpl_710 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1,
      {and_dcpl_707 , and_dcpl_710 , and_dcpl_711 , and_dcpl_714});
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      = weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      = weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_125_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = (pe_manager_base_weight_sva_mx2[14:4])
      + PEManager_15U_GetWeightAddr_else_acc_3_1;
  assign PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1[10:0];
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      = MUX_s_1_2_2(operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1, operator_3_false_1_operator_3_false_1_or_mdf_1_sva_1,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign operator_3_false_1_operator_3_false_1_or_mdf_1_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp
      = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1 | (weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1 | (weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 | (weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1) & and_dcpl_718;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 & and_dcpl_718;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1) & and_dcpl_719;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 & and_dcpl_719;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_44_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1) & and_dcpl_722;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 & and_dcpl_722;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]),
      {weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_44_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1,
      operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1, {weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse
      , and_dcpl_718 , and_dcpl_719 , and_dcpl_722});
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse
      = weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_cse,
      weight_mem_read_arbxbar_xbar_1_for_3_4_operator_7_false_1_operator_7_false_1_or_tmp);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_7_false_1_operator_7_false_1_or_tmp
      = weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1 | (weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp
      = weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_6_operator_7_false_1_operator_7_false_1_or_tmp);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_7_false_1_operator_7_false_1_or_tmp
      = Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 | (weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]));
  assign operator_7_false_1_operator_7_false_1_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 | (weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]));
  assign weight_read_addrs_0_3_0_lpi_1_dfm_4 = MUX_v_4_2_2(4'b0000, pe_manager_base_weight_sva_mx1_3_0,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_4_false_acc_sdt_sva_1 = conv_u2s_4_5(pe_config_num_manager_sva)
      + 5'b11111;
  assign operator_4_false_acc_sdt_sva_1 = nl_operator_4_false_acc_sdt_sva_1[4:0];
  assign while_and_1148_cse_1 = (~ while_if_and_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_if_and_tmp_1 = PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      = ~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl = start_PopNB_mioi_data_rsc_z_mxwt
      & pe_config_is_valid_sva & start_PopNB_mioi_return_rsc_z_mxwt;
  assign PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl = pe_config_is_zero_first_sva
      & pe_manager_zero_active_sva;
  assign PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl = ~(pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign PECore_UpdateFSM_switch_lp_mux1h_14_nl = MUX1HOT_s_1_4_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl,
      PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl, pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1,
      PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl, {PECore_UpdateFSM_switch_lp_and_7_itm_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_2_1 , PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_5_1});
  assign PECore_UpdateFSM_next_state_0_lpi_1_dfm_4 = PECore_UpdateFSM_switch_lp_mux1h_14_nl
      & PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  assign pe_config_UpdateManagerCounter_if_if_unequal_tmp = pe_config_output_counter_sva
      != (operator_8_false_acc_sdt_sva_1[7:0]);
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      = ~(pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]));
  assign input_write_req_valid_lpi_1_dfm_5 = PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      & PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1 = ~(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign PECore_RunScale_if_for_8_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_6_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[111:96]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[111:96]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[95:80]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[79:64]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[63:48]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[47:32]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[31:16]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[15:0]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[111:96]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[95:80]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[79:64]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[63:48]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[47:32]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[31:16]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[15:0]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[63:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55 , reg_weight_mem_run_3_for_5_and_162_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_163_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2
      , reg_weight_mem_run_3_for_5_and_165_itm_2_cse , reg_weight_mem_run_3_for_5_and_166_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2 , reg_weight_mem_run_3_for_5_and_168_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[79:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[95:80]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_57
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[111:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_57
      , reg_weight_mem_run_3_for_5_and_162_itm_2_cse , reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_2 , reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_3 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_3
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_3});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_96 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[15:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[31:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_96 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[47:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000004
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[63:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000005
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[79:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_96 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000006
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[95:80]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_89_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_89_nl , weight_mem_run_3_for_5_asn_306
      , weight_mem_run_3_for_5_asn_308 , reg_weight_mem_run_3_for_5_and_20_itm_2_cse
      , weight_mem_run_3_for_5_asn_310 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , weight_mem_run_3_for_5_asn_312});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_81_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_2
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[15:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_81_nl , weight_mem_run_3_for_5_asn_306
      , weight_mem_run_3_for_5_asn_308 , reg_weight_mem_run_3_for_5_and_20_itm_2_cse
      , weight_mem_run_3_for_5_asn_310 , reg_weight_mem_run_3_for_5_and_30_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_2_cse , weight_mem_run_3_for_5_asn_312});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_73_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[31:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_73_nl , weight_mem_run_3_for_5_asn_306
      , weight_mem_run_3_for_5_asn_308 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1
      , weight_mem_run_3_for_5_asn_310 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_2 , weight_mem_run_3_for_5_asn_312});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse = reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[47:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse , weight_mem_run_3_for_5_asn_306
      , weight_mem_run_3_for_5_asn_308 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2
      , weight_mem_run_3_for_5_asn_310 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_2 , weight_mem_run_3_for_5_asn_312});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 = (weight_read_addrs_1_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 = (weight_read_addrs_1_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 = (weight_read_addrs_1_lpi_1_dfm_3_2_0==3'b100)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1 = (weight_read_addrs_1_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_8_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_5_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0,
      or_dcpl_308);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      = MUX_s_1_2_2(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0,
      or_dcpl_308);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      = MUX_s_1_2_2(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0,
      or_dcpl_308);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0
      = MUX_s_1_2_2(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0,
      or_dcpl_308);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0,
      or_dcpl_308);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0,
      or_dcpl_308);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0,
      or_dcpl_308);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0,
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0,
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0,
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_if_1_and_8_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_if_1_and_5_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1 = and_289_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  assign nl_operator_16_false_acc_sdt_sva_1 = conv_u2s_8_9(pe_manager_num_input_sva)
      + 9'b111111111;
  assign operator_16_false_acc_sdt_sva_1 = nl_operator_16_false_acc_sdt_sva_1[8:0];
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1 = ~((state_mux_1_cse!=2'b00)
      | state_0_sva_mx1);
  assign PECore_UpdateFSM_switch_lp_nor_tmp_1 = ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_6 | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1
      | PECore_RunScale_PECore_RunScale_if_and_1_svs_1 | PECore_PushOutput_PECore_PushOutput_if_and_svs_1);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_87_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[127:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_87_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_80_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_80_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_111_96_sva_1
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_39_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_nl,
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_88_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[111:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_88_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_81_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[111:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_81_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_95_80_sva_1
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_nl,
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_89_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[95:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_89_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_82_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[95:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_82_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_79_64_sva_1
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_37_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_nl,
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_90_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[79:64]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_90_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_83_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[79:64]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_83_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_63_48_sva_1
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_36_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_nl,
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3);
  assign while_and_30_tmp = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp
      = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2) | reg_rva_in_reg_rw_sva_2_cse
      | (~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp!=8'b00000000))) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7])));
  assign PECore_DecodeAxiWrite_switch_lp_or_5_cse_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  assign rva_out_reg_data_63_sva_dfm_7 = PECore_PushAxiRsp_mux_18_itm_1 & rva_in_reg_rw_sva_5;
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_1_0_sva_1 = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]!=2'b00));
  assign input_mem_banks_write_if_for_if_and_stg_1_1_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b01);
  assign input_mem_banks_write_if_for_if_and_stg_1_2_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b10);
  assign input_mem_banks_write_if_for_if_and_stg_1_3_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b11);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign nl_PEManager_15U_GetInputAddr_acc_nl = input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt
      + (pe_manager_base_input_sva[7:0]);
  assign PEManager_15U_GetInputAddr_acc_nl = nl_PEManager_15U_GetInputAddr_acc_nl[7:0];
  assign input_write_addrs_lpi_1_dfm_2 = PEManager_15U_GetInputAddr_acc_nl & ({{7{PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1}},
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1})
      & ({{7{PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1}}, PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1});
  assign input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1 = ~((input_write_addrs_lpi_1_dfm_2[1:0]!=2'b00));
  assign input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b01);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b10);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b11);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2
      | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_4 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0011);
  assign PECore_DecodeAxiRead_switch_lp_nor_13_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_not_185 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 =
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:1]!=15'b000000000000000));
  assign PECore_PushAxiRsp_if_asn_59 = (~ rva_in_reg_rw_sva_10) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_61 = rva_in_reg_rw_sva_10 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_63 = input_read_req_valid_lpi_1_dfm_1_10 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign PECore_RunMac_asn_24 = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_10)
      | PECore_RunMac_PECore_RunMac_if_and_svs_10;
  assign weight_mem_run_3_for_5_asn_290 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_292 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_294 = (weight_read_addrs_7_lpi_1_dfm_3_2_0[2])
      & nor_419_cse & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_296 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_298 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_300 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_302 = (weight_read_addrs_5_lpi_1_dfm_3_2_0[2])
      & nor_425_cse & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_304 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_306 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_308 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_310 = (weight_read_addrs_3_lpi_1_dfm_3_2_0[2])
      & nor_428_cse & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_312 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign while_asn_631 = while_if_and_tmp_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign PECore_RunMac_or_cse = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_9)
      | PECore_RunMac_PECore_RunMac_if_and_svs_9;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[2:1]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_35 = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign while_and_29_cse = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign PECore_PushAxiRsp_if_asn_67 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign PECore_PushAxiRsp_if_asn_69 = (~ rva_in_reg_rw_sva_5) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign PECore_PushAxiRsp_if_asn_71 = rva_in_reg_rw_sva_5 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_96 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_166 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_168 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_7_itm_1
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_172 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_174 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_2
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_57 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_3
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_28 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_1_tmp
      = MUX_s_1_2_2(nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_3_mux_mx0w1,
      nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_mx0w0,
      operator_3_false_1_operator_3_false_1_or_mdf_1_sva_1);
  assign nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_tmp
      = MUX_s_1_2_2(operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1,
      operator_4_false_2_operator_4_false_2_or_mdf_1_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_mux_583_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1331_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_583_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_584_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1330_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_584_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_585_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1329_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_585_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_586_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1328_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_586_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_587_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1327_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_587_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_588_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1326_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_588_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1325_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_589_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1324_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_589_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_590_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1323_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_590_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_591_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1322_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_591_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_592_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1321_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_592_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_593_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1320_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_593_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_594_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1319_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_594_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1318_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1283_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_dcpl_6 = while_stage_0_11 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9;
  assign and_dcpl_7 = and_dcpl_6 & (~ rva_in_reg_rw_sva_st_1_9);
  assign and_dcpl_10 = ~(input_read_req_valid_lpi_1_dfm_1_9 | rva_in_reg_rw_sva_9);
  assign and_dcpl_28 = while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9);
  assign and_dcpl_35 = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8);
  assign and_dcpl_41 = while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign and_dcpl_45 = while_stage_0_8 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6);
  assign and_dcpl_48 = while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_11_nl = rva_in_reg_rw_sva_st_1_5 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_730_nl = rva_in_reg_rw_sva_st_1_5 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign mux_tmp = MUX_s_1_2_2(or_11_nl, and_730_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_5);
  assign mux_2_itm = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_dcpl_59 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign and_dcpl_71 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_dcpl_78 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_80 = (((Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1) | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1)
      & and_dcpl_78;
  assign and_dcpl_82 = weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign or_dcpl_28 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1;
  assign or_dcpl_31 = ((or_dcpl_28 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1) | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  assign and_dcpl_84 = or_dcpl_31 & and_dcpl_78;
  assign and_dcpl_86 = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign or_dcpl_35 = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse;
  assign and_dcpl_88 = (((Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 | or_dcpl_35) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1)
      | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp)
      & and_dcpl_78;
  assign or_dcpl_42 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse;
  assign and_dcpl_90 = (((or_dcpl_42 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1) | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1)
      & and_dcpl_78;
  assign or_dcpl_52 = ((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1) | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
  assign and_dcpl_92 = or_dcpl_52 & and_dcpl_78;
  assign or_dcpl_53 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse;
  assign or_dcpl_59 = ((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse | or_dcpl_53
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1)
      | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  assign and_dcpl_94 = or_dcpl_59 & and_dcpl_78;
  assign or_dcpl_60 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4);
  assign nor_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]));
  assign nor_197_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]));
  assign nor_198_cse = ~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]));
  assign nor_199_cse = ~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]));
  assign nor_200_cse = ~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]));
  assign and_108_cse = nor_200_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]))) & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])));
  assign nor_204_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]));
  assign and_115_cse = nor_204_cse & (~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])));
  assign or_dcpl_63 = and_115_cse | or_dcpl_60;
  assign nor_208_cse = ~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]));
  assign and_122_cse = nor_208_cse & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])));
  assign or_dcpl_64 = and_122_cse | or_dcpl_60;
  assign and_129_cse = (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) |
      (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2])));
  assign nor_218_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]));
  assign nor_219_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]));
  assign nor_216_cse = ~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]));
  assign nor_217_cse = ~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]));
  assign and_dcpl_136 = nor_216_cse & nor_217_cse & nor_218_cse & nor_219_cse;
  assign and_dcpl_137 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign and_dcpl_138 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign and_dcpl_139 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]));
  assign and_dcpl_140 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]));
  assign and_dcpl_141 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]));
  assign and_dcpl_142 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign and_dcpl_143 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign and_dcpl_144 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign and_dcpl_146 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_154 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign or_103_nl = and_741_cse | and_dcpl_136;
  assign or_100_nl = and_742_cse | and_dcpl_136;
  assign mux_tmp_13 = MUX_s_1_2_2(or_103_nl, or_100_nl, nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_tmp);
  assign and_733_cse = ((~(weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp))
      | nvhls_leading_ones_7U_nvhls_nvhls_t_7U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_1_tmp
      | Arbiter_8U_Roundrobin_pick_1_if_1_and_8_tmp | Arbiter_8U_Roundrobin_pick_1_if_1_and_5_tmp)
      & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
  assign or_tmp_27 = and_733_cse | and_dcpl_136;
  assign or_tmp_28 = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp
      | and_dcpl_136;
  assign mux_tmp_14 = MUX_s_1_2_2(or_tmp_28, or_tmp_27, weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_734_cse = Arbiter_8U_Roundrobin_pick_1_if_1_and_8_tmp | Arbiter_8U_Roundrobin_pick_1_if_1_and_5_tmp;
  assign or_110_nl = and_734_cse | and_dcpl_136;
  assign mux_tmp_15 = MUX_s_1_2_2(or_110_nl, or_tmp_27, weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign mux_tmp_16 = MUX_s_1_2_2(mux_tmp_15, mux_tmp_14, nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_tmp);
  assign or_111_cse = (~ nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_tmp)
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign mux_tmp_18 = MUX_s_1_2_2(mux_tmp_15, mux_tmp_14, or_111_cse);
  assign mux_372_nl = MUX_s_1_2_2(or_tmp_28, or_tmp_27, weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign mux_20_nl = MUX_s_1_2_2(or_tmp_28, mux_372_nl, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign mux_19_nl = MUX_s_1_2_2(or_tmp_28, or_tmp_27, and_740_cse);
  assign mux_21_nl = MUX_s_1_2_2(mux_20_nl, mux_19_nl, Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7);
  assign mux_22_nl = MUX_s_1_2_2(mux_21_nl, mux_tmp_18, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]);
  assign mux_23_nl = MUX_s_1_2_2(mux_22_nl, mux_tmp_14, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign mux_24_nl = MUX_s_1_2_2(mux_23_nl, mux_tmp_18, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign mux_25_nl = MUX_s_1_2_2(mux_24_nl, mux_tmp_14, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign mux_26_nl = MUX_s_1_2_2(mux_25_nl, mux_tmp_16, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign mux_tmp_27 = MUX_s_1_2_2(mux_26_nl, mux_tmp_14, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign and_dcpl_167 = and_dcpl_146 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]);
  assign and_dcpl_168 = and_dcpl_146 & and_dcpl_140;
  assign and_dcpl_169 = and_dcpl_146 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]);
  assign and_dcpl_170 = and_dcpl_146 & and_dcpl_139;
  assign and_dcpl_172 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_173 = and_dcpl_142 & and_dcpl_146;
  assign and_dcpl_175 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_176 = and_dcpl_141 & and_dcpl_146;
  assign and_dcpl_177 = and_dcpl_146 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]);
  assign and_dcpl_178 = and_dcpl_146 & and_dcpl_137;
  assign and_dcpl_179 = and_dcpl_146 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]);
  assign and_dcpl_180 = and_dcpl_146 & and_dcpl_138;
  assign and_dcpl_182 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_183 = and_dcpl_144 & and_dcpl_146;
  assign and_dcpl_185 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_186 = and_dcpl_143 & and_dcpl_146;
  assign and_dcpl_189 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign and_dcpl_193 = (state_2_1_sva==2'b01) & (~ state_0_sva) & and_628_cse;
  assign mux_32_nl = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      state_2_1_sva[1]);
  assign and_736_nl = (state_2_1_sva[1]) & PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  assign mux_33_nl = MUX_s_1_2_2(mux_32_nl, and_736_nl, state_2_1_sva[0]);
  assign mux_34_nl = MUX_s_1_2_2(mux_33_nl, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      state_0_sva);
  assign and_dcpl_196 = mux_34_nl & (~(PECore_RunFSM_switch_lp_nor_tmp_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign and_dcpl_197 = rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign or_dcpl_132 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]!=2'b01);
  assign and_dcpl_203 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01);
  assign and_dcpl_204 = and_dcpl_203 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]))
      & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign and_dcpl_207 = and_dcpl_204 & reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_208 = reg_rva_in_PopNB_mioi_iswt0_cse & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_210 = and_dcpl_204 & and_dcpl_208 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_212 = while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign and_dcpl_216 = weight_mem_run_3_for_land_3_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign and_dcpl_220 = weight_mem_run_3_for_land_7_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign mux_tmp_41 = MUX_s_1_2_2(and_734_cse, and_733_cse, weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign mux_tmp_42 = MUX_s_1_2_2(mux_tmp_41, mux_256_cse, nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_tmp);
  assign mux_tmp_44 = MUX_s_1_2_2(mux_tmp_41, mux_256_cse, or_111_cse);
  assign and_dcpl_237 = while_stage_0_10 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8;
  assign and_dcpl_238 = and_dcpl_197 & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_241 = and_dcpl_237 & (~ rva_in_reg_rw_sva_st_1_8);
  assign and_dcpl_252 = and_dcpl_241 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6
      | rva_in_reg_rw_sva_8 | input_read_req_valid_lpi_1_dfm_1_8));
  assign or_tmp_54 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 |
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 | rva_in_reg_rw_sva_4
      | rva_in_reg_rw_sva_st_1_4;
  assign not_tmp_147 = ~(rva_in_reg_rw_sva_4 | rva_in_reg_rw_sva_st_1_4);
  assign or_205_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      | not_tmp_147;
  assign mux_tmp_56 = MUX_s_1_2_2(or_205_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1);
  assign and_dcpl_265 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign and_dcpl_266 = and_dcpl_265 & while_stage_0_6;
  assign or_tmp_59 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      | (~ and_dcpl_212);
  assign or_tmp_60 = weight_mem_run_3_for_land_1_lpi_1_dfm_2 | (~ and_dcpl_212);
  assign mux_64_nl = MUX_s_1_2_2(or_tmp_60, or_tmp_59, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_tmp_65 = MUX_s_1_2_2((~ and_dcpl_212), mux_64_nl, while_stage_0_6);
  assign or_tmp_61 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      | and_dcpl_212;
  assign mux_66_nl = MUX_s_1_2_2((~ or_tmp_60), or_tmp_61, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_tmp_67 = MUX_s_1_2_2(and_dcpl_212, mux_66_nl, while_stage_0_6);
  assign or_tmp_63 = (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign or_215_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign mux_73_nl = MUX_s_1_2_2(or_215_nl, or_tmp_63, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_213_nl = weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign mux_74_nl = MUX_s_1_2_2(mux_73_nl, or_213_nl, weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_tmp_75 = MUX_s_1_2_2(mux_74_nl, or_tmp_63, weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_tmp_67 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | mux_tmp_75;
  assign mux_tmp_76 = MUX_s_1_2_2((~ mux_tmp_75), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_dcpl_279 = PECore_RunFSM_switch_lp_equal_tmp_1_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_292 = and_dcpl_203 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]))
      & and_dcpl_197;
  assign and_dcpl_297 = while_stage_0_9 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  assign and_dcpl_325 = and_dcpl_297 & (~ rva_in_reg_rw_sva_st_1_7);
  assign and_dcpl_354 = and_dcpl_325 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5
      | input_read_req_valid_lpi_1_dfm_1_7 | rva_in_reg_rw_sva_7));
  assign and_dcpl_362 = while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  assign and_dcpl_365 = ~(rva_in_reg_rw_sva_st_1_6 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4);
  assign and_dcpl_379 = and_dcpl_365 & (~ rva_in_reg_rw_sva_6);
  assign and_dcpl_393 = and_dcpl_212 & (~ rva_in_reg_rw_sva_st_1_5);
  assign and_dcpl_400 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | rva_in_reg_rw_sva_5);
  assign and_dcpl_438 = ~(pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1);
  assign and_dcpl_443 = and_dcpl_438 & (~ input_read_req_valid_lpi_1_dfm_1_3);
  assign or_dcpl_198 = (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp)
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp;
  assign and_dcpl_461 = or_dcpl_198 & (~(reg_rva_in_reg_rw_sva_2_cse | input_read_req_valid_lpi_1_dfm_1_2));
  assign and_dcpl_468 = or_dcpl_198 & (~ reg_rva_in_reg_rw_sva_2_cse);
  assign and_dcpl_481 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | input_read_req_valid_lpi_1_dfm_1_1);
  assign and_dcpl_482 = and_dcpl_481 & and_dcpl_189;
  assign mux_tmp_92 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1!=4'b0100));
  assign and_dcpl_488 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1);
  assign nand_17_cse = ~(PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]));
  assign and_dcpl_523 = PECore_RunMac_PECore_RunMac_if_and_svs_st_6 & while_stage_0_8
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6);
  assign and_dcpl_527 = while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
  assign or_tmp_79 = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8) | PECore_RunMac_PECore_RunMac_if_and_svs_8
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8
      | (~ while_stage_0_10);
  assign and_dcpl_536 = and_dcpl_71 & (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign nor_tmp_17 = weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & while_stage_0_7;
  assign nor_285_nl = ~(weight_mem_run_3_for_5_and_28_itm_1 | (~(weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
      & while_stage_0_7)));
  assign not_tmp_249 = MUX_s_1_2_2(nor_tmp_17, nor_285_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_dcpl_538 = and_dcpl_71 & (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign and_746_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & while_stage_0_7;
  assign nor_286_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3)
      | weight_mem_run_3_for_5_and_22_itm_1 | (~ while_stage_0_7));
  assign not_tmp_252 = MUX_s_1_2_2(and_746_nl, nor_286_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_304_nl = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  assign mux_tmp_102 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1,
      or_304_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_303_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign mux_103_nl = MUX_s_1_2_2(mux_tmp_102, or_303_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp = while_stage_0_5 & mux_103_nl;
  assign or_308_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign mux_106_nl = MUX_s_1_2_2(or_dcpl_52, or_308_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_1 = while_stage_0_5 & mux_106_nl;
  assign or_tmp_105 = Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 | and_739_cse;
  assign or_315_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign mux_109_nl = MUX_s_1_2_2(or_tmp_105, or_315_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_2 = while_stage_0_5 & mux_109_nl;
  assign or_tmp_109 = ((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1)
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  assign or_320_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_3 | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign mux_112_nl = MUX_s_1_2_2(or_tmp_109, or_320_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_3 = while_stage_0_5 & mux_112_nl;
  assign or_326_nl = PECore_RunMac_PECore_RunMac_if_and_svs_st_3 | PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
  assign mux_115_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_326_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_4 = while_stage_0_5 & mux_115_nl;
  assign or_331_nl = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  assign mux_tmp_118 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1,
      or_331_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign or_330_nl = PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 | PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign mux_119_nl = MUX_s_1_2_2(mux_tmp_118, or_330_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_5 = while_stage_0_5 & mux_119_nl;
  assign or_tmp_121 = pe_manager_zero_active_sva & pe_config_is_zero_first_sva &
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1;
  assign and_751_cse = pe_config_is_valid_sva & PECore_UpdateFSM_switch_lp_and_7_itm_1;
  assign nand_tmp_1 = ~(pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
      & (~(and_751_cse | or_tmp_121)));
  assign or_tmp_123 = and_751_cse | or_tmp_121;
  assign or_tmp_129 = state_0_sva | (state_2_1_sva!=2'b00);
  assign and_dcpl_561 = (~ weight_mem_run_3_for_land_3_lpi_1_dfm_3) & fsm_output;
  assign or_dcpl_219 = (~ while_stage_0_8) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  assign or_dcpl_222 = (~ while_stage_0_7) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign and_dcpl_579 = nor_cse & nor_197_cse;
  assign and_dcpl_580 = and_dcpl_579 & nor_198_cse & nor_199_cse;
  assign and_dcpl_582 = (~(while_stage_0_4 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
      & while_stage_0_5;
  assign or_dcpl_225 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ while_stage_0_5);
  assign and_dcpl_614 = nor_218_cse & nor_219_cse;
  assign and_dcpl_618 = nor_216_cse & nor_217_cse & and_dcpl_614;
  assign or_dcpl_226 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ while_stage_0_3);
  assign or_dcpl_231 = nand_58_cse | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_233 = or_dcpl_132 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]);
  assign and_dcpl_625 = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) |
      (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]));
  assign and_dcpl_636 = ~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]) |
      (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]));
  assign or_dcpl_273 = (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | nand_17_cse;
  assign and_dcpl_639 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]));
  assign and_dcpl_643 = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2:1]==2'b10);
  assign or_dcpl_277 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6);
  assign and_dcpl_652 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]));
  assign and_dcpl_655 = ~(weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_dcpl_665 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign and_dcpl_666 = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign or_dcpl_279 = rva_in_reg_rw_sva_6 | (~ while_stage_0_8) | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6);
  assign nor_tmp_38 = while_mux_1327_tmp & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign or_tmp_138 = ((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) & while_mux_1326_tmp)
      | nor_tmp_38;
  assign or_tmp_139 = ((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]) & while_mux_1325_tmp)
      | or_tmp_138;
  assign nor_tmp_41 = weight_mem_read_arbxbar_arbiters_next_7_5_sva & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign or_tmp_140 = ((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_6_sva)
      | nor_tmp_41;
  assign or_tmp_141 = ((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1)
      | or_tmp_140;
  assign mux_tmp_137 = MUX_s_1_2_2(or_tmp_141, or_tmp_139, while_stage_0_5);
  assign nand_3_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      & (~ or_tmp_141));
  assign mux_141_nl = MUX_s_1_2_2(nand_3_nl, or_tmp_141, and_882_cse);
  assign mux_142_nl = MUX_s_1_2_2(mux_141_nl, or_tmp_141, and_881_cse);
  assign mux_143_nl = MUX_s_1_2_2(mux_142_nl, or_tmp_141, and_880_cse);
  assign nand_2_nl = ~(while_mux_1328_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      & (~ or_tmp_139));
  assign mux_138_nl = MUX_s_1_2_2(nand_2_nl, or_tmp_139, and_886_cse);
  assign mux_139_nl = MUX_s_1_2_2(mux_138_nl, or_tmp_139, and_885_cse);
  assign mux_140_nl = MUX_s_1_2_2(mux_139_nl, or_tmp_139, and_884_cse);
  assign mux_144_itm = MUX_s_1_2_2(mux_143_nl, mux_140_nl, while_stage_0_5);
  assign or_tmp_144 = (~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])) |
      (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign mux_148_nl = MUX_s_1_2_2(nor_cse, or_tmp_144, weight_mem_read_arbxbar_arbiters_next_7_5_sva);
  assign or_435_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva | nor_tmp_41;
  assign mux_149_nl = MUX_s_1_2_2(mux_148_nl, or_435_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign or_434_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | or_tmp_140;
  assign mux_150_nl = MUX_s_1_2_2(mux_149_nl, or_434_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign nor_326_nl = ~(and_880_cse | and_881_cse | and_882_cse | and_883_cse | mux_150_nl);
  assign mux_145_nl = MUX_s_1_2_2(nor_cse, or_tmp_144, while_mux_1327_tmp);
  assign or_428_nl = while_mux_1326_tmp | nor_tmp_38;
  assign mux_146_nl = MUX_s_1_2_2(mux_145_nl, or_428_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign or_427_nl = while_mux_1325_tmp | or_tmp_138;
  assign mux_147_nl = MUX_s_1_2_2(mux_146_nl, or_427_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign nor_327_nl = ~(and_884_cse | and_885_cse | and_886_cse | and_887_cse | mux_147_nl);
  assign not_tmp_388 = MUX_s_1_2_2(nor_326_nl, nor_327_nl, while_stage_0_5);
  assign or_tmp_155 = and_886_cse | and_887_cse;
  assign or_tmp_161 = and_882_cse | and_883_cse;
  assign nor_328_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])));
  assign nor_329_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_3_sva | and_883_cse);
  assign mux_155_nl = MUX_s_1_2_2(nor_328_nl, nor_329_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nor_330_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_1_sva | or_tmp_161);
  assign mux_156_nl = MUX_s_1_2_2(mux_155_nl, nor_330_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign nor_331_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_2_sva | and_881_cse
      | or_tmp_161);
  assign mux_157_nl = MUX_s_1_2_2(mux_156_nl, nor_331_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign nor_332_nl = ~(while_mux_1328_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])));
  assign nor_333_nl = ~(while_mux_1329_tmp | and_887_cse);
  assign mux_152_nl = MUX_s_1_2_2(nor_332_nl, nor_333_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nor_334_nl = ~(while_mux_1331_tmp | or_tmp_155);
  assign mux_153_nl = MUX_s_1_2_2(mux_152_nl, nor_334_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign nor_335_nl = ~(while_mux_1330_tmp | and_885_cse | or_tmp_155);
  assign mux_154_nl = MUX_s_1_2_2(mux_153_nl, nor_335_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign mux_158_nl = MUX_s_1_2_2(mux_157_nl, mux_154_nl, while_stage_0_5);
  assign and_dcpl_674 = mux_158_nl & and_dcpl_579;
  assign and_782_cse = while_mux_1318_tmp & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_tmp_175 = ((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & while_mux_1320_tmp)
      | and_782_cse;
  assign or_tmp_177 = ((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_5_sva)
      | (Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]));
  assign or_463_nl = and_888_cse | or_tmp_177;
  assign or_461_nl = and_893_cse | or_tmp_175;
  assign mux_tmp_160 = MUX_s_1_2_2(or_463_nl, or_461_nl, while_stage_0_5);
  assign nand_5_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      & (~ or_tmp_177));
  assign mux_164_nl = MUX_s_1_2_2(nand_5_nl, or_tmp_177, and_891_cse);
  assign mux_165_nl = MUX_s_1_2_2(mux_164_nl, or_tmp_177, and_890_cse);
  assign mux_166_nl = MUX_s_1_2_2(mux_165_nl, or_tmp_177, and_889_cse);
  assign nor_336_nl = ~(and_888_cse | mux_166_nl);
  assign nand_4_nl = ~(while_mux_1324_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      & (~ or_tmp_175));
  assign mux_161_nl = MUX_s_1_2_2(nand_4_nl, or_tmp_175, and_896_cse);
  assign mux_162_nl = MUX_s_1_2_2(mux_161_nl, or_tmp_175, and_895_cse);
  assign mux_163_nl = MUX_s_1_2_2(mux_162_nl, or_tmp_175, and_894_cse);
  assign nor_337_nl = ~(and_893_cse | mux_163_nl);
  assign not_tmp_393 = MUX_s_1_2_2(nor_336_nl, nor_337_nl, while_stage_0_5);
  assign or_tmp_182 = and_782_cse | and_893_cse;
  assign or_470_nl = while_mux_1319_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign or_469_nl = while_mux_1318_tmp | and_893_cse;
  assign mux_168_nl = MUX_s_1_2_2(or_470_nl, or_469_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_169_nl = MUX_s_1_2_2(mux_168_nl, or_tmp_182, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_468_nl = while_mux_1320_tmp | or_tmp_182;
  assign mux_170_nl = MUX_s_1_2_2(mux_169_nl, or_468_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_187 = and_896_cse | and_895_cse | mux_170_nl;
  assign or_tmp_190 = and_888_cse | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  assign mux_tmp_171 = MUX_s_1_2_2(and_888_cse, or_tmp_190, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_477_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign mux_172_nl = MUX_s_1_2_2(or_477_nl, or_tmp_190, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_173_nl = MUX_s_1_2_2(mux_172_nl, mux_tmp_171, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_476_nl = weight_mem_read_arbxbar_arbiters_next_6_5_sva | mux_tmp_171;
  assign mux_174_nl = MUX_s_1_2_2(mux_173_nl, or_476_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_194 = and_891_cse | and_890_cse | mux_174_nl;
  assign mux_179_nl = MUX_s_1_2_2(or_tmp_194, or_tmp_187, while_stage_0_5);
  assign or_484_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | or_tmp_194;
  assign or_483_nl = while_mux_1322_tmp | or_tmp_187;
  assign mux_178_nl = MUX_s_1_2_2(or_484_nl, or_483_nl, while_stage_0_5);
  assign mux_180_nl = MUX_s_1_2_2(mux_179_nl, mux_178_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign or_482_nl = weight_mem_read_arbxbar_arbiters_next_6_1_sva | or_tmp_194;
  assign or_481_nl = while_mux_1324_tmp | or_tmp_187;
  assign mux_176_nl = MUX_s_1_2_2(or_482_nl, or_481_nl, while_stage_0_5);
  assign or_480_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | or_tmp_194;
  assign or_473_nl = while_mux_1322_tmp | while_mux_1324_tmp | or_tmp_187;
  assign mux_175_nl = MUX_s_1_2_2(or_480_nl, or_473_nl, while_stage_0_5);
  assign mux_177_nl = MUX_s_1_2_2(mux_176_nl, mux_175_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_181_itm = MUX_s_1_2_2(mux_180_nl, mux_177_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_tmp_200 = and_896_cse | and_897_cse;
  assign or_tmp_206 = and_891_cse | and_892_cse;
  assign nor_338_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_1_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])));
  assign nor_339_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_2_sva | and_892_cse);
  assign mux_185_nl = MUX_s_1_2_2(nor_338_nl, nor_339_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign nor_340_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_4_sva | or_tmp_206);
  assign mux_186_nl = MUX_s_1_2_2(mux_185_nl, nor_340_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign nor_341_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_3_sva | and_890_cse
      | or_tmp_206);
  assign mux_187_nl = MUX_s_1_2_2(mux_186_nl, nor_341_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nor_342_nl = ~(while_mux_1324_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])));
  assign nor_343_nl = ~(while_mux_1323_tmp | and_897_cse);
  assign mux_182_nl = MUX_s_1_2_2(nor_342_nl, nor_343_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign nor_344_nl = ~(while_mux_1321_tmp | or_tmp_200);
  assign mux_183_nl = MUX_s_1_2_2(mux_182_nl, nor_344_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign nor_345_nl = ~(while_mux_1322_tmp | and_895_cse | or_tmp_200);
  assign mux_184_nl = MUX_s_1_2_2(mux_183_nl, nor_345_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_188_nl = MUX_s_1_2_2(mux_187_nl, mux_184_nl, while_stage_0_5);
  assign and_dcpl_677 = mux_188_nl & nor_200_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])));
  assign nor_tmp_116 = weight_mem_read_arbxbar_arbiters_next_5_5_sva & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign and_812_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1;
  assign or_510_nl = and_812_cse | nor_tmp_116;
  assign and_814_nl = Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign mux_190_nl = MUX_s_1_2_2(nor_tmp_116, and_814_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_509_nl = ((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]) & Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1)
      | mux_190_nl;
  assign or_508_nl = and_812_cse | (Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_cse
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]));
  assign mux_191_nl = MUX_s_1_2_2(or_509_nl, or_508_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_192 = MUX_s_1_2_2(or_510_nl, mux_191_nl, while_stage_0_5);
  assign and_dcpl_678 = mux_tmp_192 | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  assign and_dcpl_680 = (~ mux_tmp_192) & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp)
      & weight_mem_read_arbxbar_xbar_1_for_3_6_operator_7_false_1_operator_7_false_1_or_tmp;
  assign and_dcpl_681 = ~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]))) | weight_mem_read_arbxbar_xbar_1_for_3_6_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_dcpl_684 = nor_204_cse & (~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]))
      & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]) | weight_mem_read_arbxbar_xbar_1_for_3_6_operator_7_false_1_operator_7_false_1_or_tmp));
  assign Arbiter_8U_Roundrobin_pick_1_mux_605_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign mux_194_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_605_nl, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_cse,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_195 = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_5_sva,
      mux_194_nl, while_stage_0_5);
  assign and_dcpl_686 = (mux_tmp_195 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]))
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  assign and_dcpl_689 = (~(mux_tmp_195 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])))
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp))
      & weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp;
  assign and_dcpl_690 = ~((~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]))) | weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_dcpl_693 = nor_208_cse & (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]))
      & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]) | weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp));
  assign and_dcpl_695 = ~(weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp);
  assign nor_tmp_121 = weight_mem_read_arbxbar_arbiters_next_2_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign or_tmp_228 = ((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_3_sva)
      | nor_tmp_121;
  assign or_tmp_229 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_1_sva)
      | or_tmp_228;
  assign or_tmp_230 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_2_sva)
      | or_tmp_229;
  assign nor_tmp_125 = Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign or_tmp_231 = ((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]) & Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1)
      | nor_tmp_125;
  assign or_tmp_232 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]) & Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1)
      | or_tmp_231;
  assign or_530_nl = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) & Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1)
      | or_tmp_232;
  assign mux_197_nl = MUX_s_1_2_2(or_tmp_230, or_530_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_524_nl = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign mux_196_nl = MUX_s_1_2_2(or_tmp_230, or_524_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign mux_198_nl = MUX_s_1_2_2(mux_197_nl, mux_196_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_199 = MUX_s_1_2_2(or_tmp_230, mux_198_nl, while_stage_0_5);
  assign and_dcpl_696 = mux_tmp_199 & and_dcpl_695;
  assign and_dcpl_697 = (~((~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]))) | mux_tmp_199)) &
      and_dcpl_695;
  assign or_535_nl = weight_mem_read_arbxbar_arbiters_next_2_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]));
  assign or_534_nl = weight_mem_read_arbxbar_arbiters_next_2_3_sva | nor_tmp_121;
  assign mux_200_nl = MUX_s_1_2_2(or_535_nl, or_534_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign or_533_nl = weight_mem_read_arbxbar_arbiters_next_2_1_sva | or_tmp_228;
  assign mux_201_nl = MUX_s_1_2_2(mux_200_nl, or_533_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign or_532_nl = weight_mem_read_arbxbar_arbiters_next_2_2_sva | or_tmp_229;
  assign mux_tmp_202 = MUX_s_1_2_2(mux_201_nl, or_532_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign or_540_nl = Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]));
  assign or_539_nl = Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 | nor_tmp_125;
  assign mux_203_nl = MUX_s_1_2_2(or_540_nl, or_539_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign or_538_nl = Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 | or_tmp_231;
  assign mux_204_nl = MUX_s_1_2_2(mux_203_nl, or_538_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign or_537_nl = Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 | or_tmp_232;
  assign mux_205_nl = MUX_s_1_2_2(mux_204_nl, or_537_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign mux_206_nl = MUX_s_1_2_2(mux_tmp_202, mux_205_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_536_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2])
      | mux_tmp_202;
  assign mux_207_nl = MUX_s_1_2_2(mux_206_nl, or_536_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_208_nl = MUX_s_1_2_2(mux_tmp_202, mux_207_nl, while_stage_0_5);
  assign and_dcpl_703 = ~(mux_208_nl | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]));
  assign nor_tmp_127 = while_mux_1283_tmp & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign or_tmp_245 = and_903_cse | nor_tmp_127;
  assign or_tmp_247 = and_910_cse | nor_tmp_127;
  assign or_tmp_250 = and_903_cse | and_904_cse;
  assign mux_212_nl = MUX_s_1_2_2(or_tmp_245, or_tmp_247, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_550_nl = (Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_cse
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])) | nor_tmp_127;
  assign mux_213_nl = MUX_s_1_2_2(mux_212_nl, or_550_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_214_nl = MUX_s_1_2_2(or_tmp_250, mux_213_nl, while_stage_0_5);
  assign or_548_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_250;
  assign or_546_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_245;
  assign or_545_nl = Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 | or_tmp_247;
  assign mux_209_nl = MUX_s_1_2_2(or_546_nl, or_545_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_543_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1])
      | weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_245;
  assign mux_210_nl = MUX_s_1_2_2(mux_209_nl, or_543_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_211_nl = MUX_s_1_2_2(or_548_nl, mux_210_nl, while_stage_0_5);
  assign mux_tmp_215 = MUX_s_1_2_2(mux_214_nl, mux_211_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign nand_7_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      & (~ or_tmp_245));
  assign mux_216_nl = MUX_s_1_2_2(nand_7_nl, or_tmp_245, and_901_cse);
  assign mux_217_nl = MUX_s_1_2_2(mux_216_nl, or_tmp_245, and_900_cse);
  assign mux_218_nl = MUX_s_1_2_2(mux_217_nl, or_tmp_245, and_898_cse);
  assign or_tmp_259 = and_899_cse | mux_218_nl;
  assign nand_9_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      & (~ or_tmp_250));
  assign mux_225_nl = MUX_s_1_2_2(nand_9_nl, or_tmp_250, and_901_cse);
  assign mux_226_nl = MUX_s_1_2_2(mux_225_nl, or_tmp_250, and_900_cse);
  assign mux_227_nl = MUX_s_1_2_2(mux_226_nl, or_tmp_250, and_898_cse);
  assign or_560_nl = and_899_cse | mux_227_nl;
  assign nand_8_nl = ~(Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      & (~ or_tmp_247));
  assign mux_220_nl = MUX_s_1_2_2(nand_8_nl, or_tmp_247, and_908_cse);
  assign mux_221_nl = MUX_s_1_2_2(mux_220_nl, or_tmp_247, and_907_cse);
  assign mux_222_nl = MUX_s_1_2_2(mux_221_nl, or_tmp_247, and_905_cse);
  assign or_558_nl = and_906_cse | mux_222_nl;
  assign mux_223_nl = MUX_s_1_2_2(or_tmp_259, or_558_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_554_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]))) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])
      | nor_tmp_127;
  assign mux_219_nl = MUX_s_1_2_2(or_tmp_259, or_554_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign mux_224_nl = MUX_s_1_2_2(mux_223_nl, mux_219_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_228_itm = MUX_s_1_2_2(or_560_nl, mux_224_nl, while_stage_0_5);
  assign or_tmp_267 = and_898_cse | and_900_cse | and_901_cse | and_902_cse;
  assign or_tmp_268 = and_903_cse | or_tmp_267;
  assign or_tmp_269 = and_899_cse | or_tmp_268;
  assign or_tmp_272 = and_905_cse | and_907_cse | and_908_cse | and_909_cse;
  assign or_tmp_273 = and_910_cse | or_tmp_272;
  assign or_577_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])) | weight_mem_read_arbxbar_arbiters_next_1_6_sva
      | or_tmp_267;
  assign mux_233_nl = MUX_s_1_2_2(or_577_nl, or_tmp_268, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign or_575_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_268;
  assign mux_tmp_234 = MUX_s_1_2_2(mux_233_nl, or_575_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign or_580_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])) | Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1
      | or_tmp_272;
  assign mux_236_nl = MUX_s_1_2_2(or_580_nl, or_tmp_273, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign or_578_nl = Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 | or_tmp_273;
  assign mux_237_nl = MUX_s_1_2_2(mux_236_nl, or_578_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign mux_238_nl = MUX_s_1_2_2(mux_tmp_234, mux_237_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_574_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | (~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]))
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign mux_235_nl = MUX_s_1_2_2(mux_tmp_234, or_574_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign mux_239_nl = MUX_s_1_2_2(mux_238_nl, mux_235_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_240_nl = MUX_s_1_2_2(mux_tmp_234, mux_239_nl, while_stage_0_5);
  assign or_573_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      | or_tmp_269;
  assign or_571_nl = and_906_cse | or_tmp_273;
  assign mux_230_nl = MUX_s_1_2_2(or_tmp_269, or_571_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_561_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign mux_229_nl = MUX_s_1_2_2(or_tmp_269, or_561_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign mux_231_nl = MUX_s_1_2_2(mux_230_nl, mux_229_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_572_nl = while_mux_1283_tmp | mux_231_nl;
  assign mux_232_nl = MUX_s_1_2_2(or_573_nl, or_572_nl, while_stage_0_5);
  assign mux_241_itm = MUX_s_1_2_2(mux_240_nl, mux_232_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign or_tmp_284 = and_898_cse | and_901_cse;
  assign or_586_nl = weight_mem_read_arbxbar_arbiters_next_1_3_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]));
  assign or_585_nl = weight_mem_read_arbxbar_arbiters_next_1_1_sva | and_901_cse;
  assign mux_242_nl = MUX_s_1_2_2(or_586_nl, or_585_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign or_584_nl = weight_mem_read_arbxbar_arbiters_next_1_2_sva | or_tmp_284;
  assign mux_243_nl = MUX_s_1_2_2(mux_242_nl, or_584_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign or_583_nl = weight_mem_read_arbxbar_arbiters_next_1_4_sva | and_900_cse
      | or_tmp_284;
  assign mux_tmp_244 = MUX_s_1_2_2(mux_243_nl, or_583_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign or_tmp_291 = and_905_cse | and_908_cse;
  assign or_593_nl = Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]));
  assign or_592_nl = Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 | and_908_cse;
  assign mux_245_nl = MUX_s_1_2_2(or_593_nl, or_592_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign or_591_nl = Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 | or_tmp_291;
  assign mux_246_nl = MUX_s_1_2_2(mux_245_nl, or_591_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign or_590_nl = Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 | and_907_cse | or_tmp_291;
  assign mux_247_nl = MUX_s_1_2_2(mux_246_nl, or_590_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign mux_248_nl = MUX_s_1_2_2(mux_tmp_244, mux_247_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign or_587_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1])
      | mux_tmp_244;
  assign mux_249_nl = MUX_s_1_2_2(mux_248_nl, or_587_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_250_nl = MUX_s_1_2_2(mux_tmp_244, mux_249_nl, while_stage_0_5);
  assign and_dcpl_705 = (~ mux_250_nl) & and_dcpl_614;
  assign or_tmp_304 = and_898_cse | and_899_cse | and_900_cse | and_901_cse | and_902_cse
      | and_903_cse | nor_tmp_127;
  assign while_mux_1335_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_255 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1,
      while_mux_1335_nl, while_stage_0_5);
  assign and_dcpl_707 = (mux_tmp_255 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]))
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  assign and_dcpl_710 = (~(mux_tmp_255 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])))
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp))
      & weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp;
  assign and_dcpl_711 = ~((~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]))) | weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_dcpl_714 = (~(weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])))
      & and_dcpl_625;
  assign and_dcpl_718 = (~(weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp))
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp)
      & weight_mem_read_arbxbar_xbar_1_for_3_4_operator_7_false_1_operator_7_false_1_or_tmp;
  assign and_dcpl_719 = ~((~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]))) | weight_mem_read_arbxbar_xbar_1_for_3_4_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_dcpl_722 = and_dcpl_636 & (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]))
      & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | weight_mem_read_arbxbar_xbar_1_for_3_4_operator_7_false_1_operator_7_false_1_or_tmp));
  assign or_dcpl_308 = ~(Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs);
  assign PECore_PushAxiRsp_mux_18_itm_1_mx0c1 = and_dcpl_212 & (~ rva_in_reg_rw_sva_5);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_a = weight_port_read_out_data_3_7_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[127:112];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_c = weight_port_read_out_data_3_6_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[111:96];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_1_a = weight_port_read_out_data_7_1_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[31:16];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_1_c = weight_port_read_out_data_7_0_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[15:0];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_2_a = weight_port_read_out_data_7_3_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[63:48];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_2_c = weight_port_read_out_data_7_2_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[47:32];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_3_a = weight_port_read_out_data_7_5_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[95:80];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_3_c = weight_port_read_out_data_7_4_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[79:64];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_4_a = weight_port_read_out_data_7_7_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_4_c = weight_port_read_out_data_7_6_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_5_a = {weight_port_read_out_data_0_1_sva_dfm_1_1_15
      , weight_port_read_out_data_0_1_sva_dfm_1_1_14_0};
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[31:16];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_5_c = {weight_port_read_out_data_0_0_sva_dfm_1_1_15
      , weight_port_read_out_data_0_0_sva_dfm_1_1_14_0};
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[15:0];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_a = {weight_port_read_out_data_0_3_sva_dfm_1_1_15
      , weight_port_read_out_data_0_3_sva_dfm_1_1_14_0};
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[63:48];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_c = {weight_port_read_out_data_0_2_sva_dfm_1_1_15
      , weight_port_read_out_data_0_2_sva_dfm_1_1_14_0};
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[47:32];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_a = weight_mem_run_3_for_5_mux_5_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[95:80];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_c = weight_mem_run_3_for_5_mux_4_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[79:64];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_8_a = weight_mem_run_3_for_5_mux_7_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[127:112];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_8_c = weight_mem_run_3_for_5_mux_6_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[111:96];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_9_a = weight_mem_run_3_for_5_mux_49_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_9_c = weight_mem_run_3_for_5_mux_48_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_10_a = weight_mem_run_3_for_5_mux_51_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_10_c = weight_mem_run_3_for_5_mux_50_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_11_a = weight_mem_run_3_for_5_mux_53_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_11_c = weight_mem_run_3_for_5_mux_52_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_12_a = weight_mem_run_3_for_5_mux_55_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_12_c = weight_mem_run_3_for_5_mux_54_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_13_a = weight_mem_run_3_for_5_mux_9_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_13_c = weight_mem_run_3_for_5_mux_8_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_14_a = rva_out_reg_data_127_112_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_14_c = rva_out_reg_data_111_96_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_15_a = rva_out_reg_data_95_80_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_15_c = rva_out_reg_data_79_64_sva_dfm_4_1;
  assign and_569_nl = fsm_output & (~ weight_mem_run_3_for_land_2_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_16_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
      weight_port_read_out_data_1_7_sva_dfm_1, and_569_nl);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_16_c = weight_mem_run_3_for_5_mux_14_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_17_a = weight_port_read_out_data_5_1_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_17_c = weight_port_read_out_data_5_0_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_18_a = weight_port_read_out_data_5_3_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_18_c = weight_port_read_out_data_5_2_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_19_a = weight_port_read_out_data_5_5_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_19_c = weight_port_read_out_data_5_4_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_20_a = weight_port_read_out_data_5_7_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_20_c = weight_port_read_out_data_5_6_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_21_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
      weight_port_read_out_data_2_1_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_21_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001,
      weight_port_read_out_data_2_0_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_22_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002,
      weight_port_read_out_data_2_3_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_22_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003,
      weight_port_read_out_data_2_2_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_23_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000004,
      weight_port_read_out_data_2_5_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_23_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000005,
      weight_port_read_out_data_2_4_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_24_a = weight_mem_run_3_for_5_mux_23_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_24_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000006,
      weight_port_read_out_data_2_6_sva_dfm_1, and_dcpl_561);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_25_a = weight_mem_run_3_for_5_mux_33_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_25_c = weight_mem_run_3_for_5_mux_32_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_26_a = weight_mem_run_3_for_5_mux_35_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_26_c = weight_mem_run_3_for_5_mux_34_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_27_a = weight_mem_run_3_for_5_mux_37_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_27_c = weight_mem_run_3_for_5_mux_36_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_28_a = weight_mem_run_3_for_5_mux_39_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_28_c = weight_mem_run_3_for_5_mux_38_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_29_a = weight_mem_run_3_for_5_mux_25_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_29_c = weight_mem_run_3_for_5_mux_24_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_30_a = weight_mem_run_3_for_5_mux_27_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_30_c = weight_mem_run_3_for_5_mux_26_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_31_a = weight_port_read_out_data_3_5_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_31_c = weight_port_read_out_data_3_4_sva_dfm_3;
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0));
  assign weight_mem_banks_write_if_for_if_and_35_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_36_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_37_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_38_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_39_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_40_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_41_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      , weight_mem_banks_write_if_for_if_and_35_nl , weight_mem_banks_write_if_for_if_and_36_nl
      , weight_mem_banks_write_if_for_if_and_37_nl , weight_mem_banks_write_if_for_if_and_38_nl
      , weight_mem_banks_write_if_for_if_and_39_nl , weight_mem_banks_write_if_for_if_and_40_nl
      , weight_mem_banks_write_if_for_if_and_41_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0});
  assign weight_mem_banks_write_if_for_if_mux_7_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      , weight_mem_banks_write_if_for_if_mux_7_nl};
  assign nor_381_nl = ~((~ PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3) |
      PECore_RunFSM_switch_lp_equal_tmp_1_2);
  assign mux_136_nl = MUX_s_1_2_2(mux_tmp_118, nor_381_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff = mux_136_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_2[14:3];
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff = and_dcpl_167;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0));
  assign weight_mem_banks_write_if_for_if_and_28_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_29_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_30_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_31_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_32_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_33_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_34_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      , weight_mem_banks_write_if_for_if_and_28_nl , weight_mem_banks_write_if_for_if_and_29_nl
      , weight_mem_banks_write_if_for_if_and_30_nl , weight_mem_banks_write_if_for_if_and_31_nl
      , weight_mem_banks_write_if_for_if_and_32_nl , weight_mem_banks_write_if_for_if_and_33_nl
      , weight_mem_banks_write_if_for_if_and_34_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0});
  assign weight_mem_banks_write_if_for_if_mux_6_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      , weight_mem_banks_write_if_for_if_mux_6_nl};
  assign nor_380_nl = ~((~ PECore_RunMac_PECore_RunMac_if_and_svs_st_3) | PECore_UpdateFSM_switch_lp_equal_tmp_2_3);
  assign mux_135_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_380_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff = mux_135_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff = and_dcpl_169;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0));
  assign weight_mem_banks_write_if_for_if_and_21_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_22_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_23_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_24_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_25_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_26_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_27_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      , weight_mem_banks_write_if_for_if_and_21_nl , weight_mem_banks_write_if_for_if_and_22_nl
      , weight_mem_banks_write_if_for_if_and_23_nl , weight_mem_banks_write_if_for_if_and_24_nl
      , weight_mem_banks_write_if_for_if_and_25_nl , weight_mem_banks_write_if_for_if_and_26_nl
      , weight_mem_banks_write_if_for_if_and_27_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0});
  assign weight_mem_banks_write_if_for_if_mux_5_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      , weight_mem_banks_write_if_for_if_mux_5_nl};
  assign nor_379_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_3) | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]));
  assign mux_134_nl = MUX_s_1_2_2(or_tmp_109, nor_379_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff = mux_134_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff = and_dcpl_172;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0));
  assign weight_mem_banks_write_if_for_if_and_14_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_15_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_16_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_17_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_18_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_19_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_20_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      , weight_mem_banks_write_if_for_if_and_14_nl , weight_mem_banks_write_if_for_if_and_15_nl
      , weight_mem_banks_write_if_for_if_and_16_nl , weight_mem_banks_write_if_for_if_and_17_nl
      , weight_mem_banks_write_if_for_if_and_18_nl , weight_mem_banks_write_if_for_if_and_19_nl
      , weight_mem_banks_write_if_for_if_and_20_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0});
  assign weight_mem_banks_write_if_for_if_mux_4_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      , weight_mem_banks_write_if_for_if_mux_4_nl};
  assign nor_378_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3) | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]));
  assign mux_133_nl = MUX_s_1_2_2(or_tmp_105, nor_378_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff = mux_133_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff = and_dcpl_175;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0));
  assign weight_mem_banks_write_if_for_if_and_7_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_9_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_10_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_11_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_12_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_13_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      , weight_mem_banks_write_if_for_if_and_7_nl , weight_mem_banks_write_if_for_if_and_8_nl
      , weight_mem_banks_write_if_for_if_and_9_nl , weight_mem_banks_write_if_for_if_and_10_nl
      , weight_mem_banks_write_if_for_if_and_11_nl , weight_mem_banks_write_if_for_if_and_12_nl
      , weight_mem_banks_write_if_for_if_and_13_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0});
  assign weight_mem_banks_write_if_for_if_mux_3_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      , weight_mem_banks_write_if_for_if_mux_3_nl};
  assign nor_377_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1)
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]));
  assign mux_132_nl = MUX_s_1_2_2(or_dcpl_52, nor_377_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff = mux_132_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff = and_dcpl_177;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0));
  assign weight_mem_banks_write_if_for_if_and_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_1_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_2_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_3_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_5_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl ,
      weight_mem_banks_write_if_for_if_and_nl , weight_mem_banks_write_if_for_if_and_1_nl
      , weight_mem_banks_write_if_for_if_and_2_nl , weight_mem_banks_write_if_for_if_and_3_nl
      , weight_mem_banks_write_if_for_if_and_4_nl , weight_mem_banks_write_if_for_if_and_5_nl
      , weight_mem_banks_write_if_for_if_and_6_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0});
  assign weight_mem_banks_write_if_for_if_mux_2_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      , weight_mem_banks_write_if_for_if_mux_2_nl};
  assign nor_376_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1)
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]));
  assign mux_131_nl = MUX_s_1_2_2(mux_tmp_102, nor_376_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff = mux_131_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff = and_dcpl_179;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_1_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_54_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0,
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_1_nl
      , weight_mem_banks_write_if_for_if_mux_54_nl};
  assign nor_375_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1);
  assign mux_130_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_375_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff = mux_130_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_3_14_3;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff = and_dcpl_538;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_53_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0,
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_nl
      , weight_mem_banks_write_if_for_if_mux_53_nl};
  assign nor_374_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_1);
  assign mux_129_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_374_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff = mux_129_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff = and_dcpl_536;
  assign and_dcpl_723 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1
      & (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign or_dcpl = and_dcpl_723 | ((weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1);
  assign and_dcpl_724 = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])
      & (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign mux_tmp_256 = MUX_s_1_2_2((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]),
      (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign or_dcpl_309 = (mux_tmp_256 & and_dcpl_639) | (and_dcpl_724 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign nor_tmp_191 = and_dcpl_265 & while_stage_0_6 & (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2])
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign or_647_cse = PECore_RunMac_PECore_RunMac_if_and_svs_9 | PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign or_dcpl_314 = ~(or_647_cse & and_dcpl_28);
  assign or_648_cse = PECore_UpdateFSM_switch_lp_equal_tmp_2_8 | PECore_RunMac_PECore_RunMac_if_and_svs_8;
  assign or_dcpl_315 = ~(or_648_cse & and_dcpl_35);
  assign or_dcpl_316 = and_dcpl_723 | ((weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1);
  assign and_647_ssc = and_dcpl_639 & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]));
  assign and_648_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign and_649_ssc = and_dcpl_639 & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign PECore_DecodeAxiRead_switch_lp_mux_21_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[0]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl
      = PECore_DecodeAxiRead_switch_lp_mux_21_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_25_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl,
      rva_out_reg_data_0_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_19_nl = MUX_s_1_2_2(rva_out_reg_data_mux_25_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_PushAxiRsp_if_mux1h_9 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_19_nl,
      (weight_port_read_out_data_0_0_sva_dfm_5_14_0[0]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl
      = (SC_SRAM_CONFIG[7:1]) & (signext_7_1(~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9))
      & ({{6{PECore_DecodeAxiRead_switch_lp_nor_9_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1});
  assign PECore_PushAxiRsp_if_mux1h_10 = MUX1HOT_v_7_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl,
      rva_out_reg_data_7_1_sva_dfm_6, input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5,
      (weight_port_read_out_data_0_0_sva_dfm_5_14_0[7:1]), {PECore_PushAxiRsp_if_asn_59
      , PECore_PushAxiRsp_if_asn_61 , PECore_PushAxiRsp_if_asn_63 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_22_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[8]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl
      = PECore_DecodeAxiRead_switch_lp_mux_22_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_26_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl,
      rva_out_reg_data_8_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_20_nl = MUX_s_1_2_2(rva_out_reg_data_mux_26_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_PushAxiRsp_if_mux1h_11 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_20_nl,
      (weight_port_read_out_data_0_0_sva_dfm_5_14_0[8]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign PECore_DecodeAxiRead_switch_lp_mux_18_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[15]),
      (rva_out_reg_data_15_9_sva_dfm_10[6]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl
      = PECore_DecodeAxiRead_switch_lp_mux_18_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_12_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl,
      rva_out_reg_data_15_9_sva_dfm_6_6, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5[6]),
      weight_port_read_out_data_0_0_sva_dfm_5_15, {PECore_PushAxiRsp_if_asn_59 ,
      PECore_PushAxiRsp_if_asn_61 , PECore_PushAxiRsp_if_asn_63 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_25_nl = MUX_v_6_2_2((SC_SRAM_CONFIG[14:9]),
      (rva_out_reg_data_15_9_sva_dfm_10[5:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl
      = MUX_v_6_2_2(6'b000000, PECore_DecodeAxiRead_switch_lp_mux_25_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_12_5_0 = MUX1HOT_v_6_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl,
      rva_out_reg_data_15_9_sva_dfm_6_5_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5[5:0]),
      (weight_port_read_out_data_0_0_sva_dfm_5_14_0[14:9]), {PECore_PushAxiRsp_if_asn_59
      , PECore_PushAxiRsp_if_asn_61 , PECore_PushAxiRsp_if_asn_63 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_23_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[16]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl
      = PECore_DecodeAxiRead_switch_lp_mux_23_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_27_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl,
      rva_out_reg_data_16_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_21_nl = MUX_s_1_2_2(rva_out_reg_data_mux_27_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_PushAxiRsp_if_mux1h_13 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_21_nl,
      (weight_port_read_out_data_0_1_sva_dfm_5_rsp_1[0]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign PECore_DecodeAxiRead_switch_lp_mux_19_nl = MUX_v_7_2_2((SC_SRAM_CONFIG[23:17]),
      rva_out_reg_data_23_17_sva_dfm_8, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl
      = MUX_v_7_2_2(7'b0000000, PECore_DecodeAxiRead_switch_lp_mux_19_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_14 = MUX1HOT_v_7_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl,
      rva_out_reg_data_23_17_sva_dfm_6, input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5,
      (weight_port_read_out_data_0_1_sva_dfm_5_rsp_1[7:1]), {PECore_PushAxiRsp_if_asn_59
      , PECore_PushAxiRsp_if_asn_61 , PECore_PushAxiRsp_if_asn_63 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_24_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[24]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl
      = PECore_DecodeAxiRead_switch_lp_mux_24_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_29_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl,
      rva_out_reg_data_24_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_22_nl = MUX_s_1_2_2(rva_out_reg_data_mux_29_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_PushAxiRsp_if_mux1h_15 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_22_nl,
      (weight_port_read_out_data_0_1_sva_dfm_5_rsp_1[8]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign PECore_DecodeAxiRead_switch_lp_mux_20_nl = MUX_v_6_2_2((SC_SRAM_CONFIG[30:25]),
      rva_out_reg_data_30_25_sva_dfm_8, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl =
      MUX_v_6_2_2(6'b000000, PECore_DecodeAxiRead_switch_lp_mux_20_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_16 = MUX1HOT_v_6_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl,
      rva_out_reg_data_30_25_sva_dfm_6, input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5,
      (weight_port_read_out_data_0_1_sva_dfm_5_rsp_1[14:9]), {PECore_PushAxiRsp_if_asn_59
      , PECore_PushAxiRsp_if_asn_61 , PECore_PushAxiRsp_if_asn_63 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl
      = (SC_SRAM_CONFIG[31]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9) &
      PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_28_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl,
      rva_out_reg_data_31_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_23_nl = MUX_s_1_2_2(rva_out_reg_data_mux_28_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_PushAxiRsp_if_mux1h_17 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_23_nl,
      weight_port_read_out_data_0_1_sva_dfm_5_rsp_0, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign nl_ProductSum_for_acc_26_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_16_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_15_z);
  assign ProductSum_for_acc_26_nl = nl_ProductSum_for_acc_26_nl[34:0];
  assign nl_ProductSum_for_acc_27_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_14_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_13_z);
  assign ProductSum_for_acc_27_nl = nl_ProductSum_for_acc_27_nl[34:0];
  assign nl_ProductSum_for_acc_25_nl = ProductSum_for_acc_26_nl + ProductSum_for_acc_27_nl;
  assign ProductSum_for_acc_25_nl = nl_ProductSum_for_acc_25_nl[34:0];
  assign PECore_UpdateFSM_switch_lp_not_37_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_1_itm
      = MUX_v_35_2_2(35'b00000000000000000000000000000000000, ProductSum_for_acc_25_nl,
      PECore_UpdateFSM_switch_lp_not_37_nl);
  assign nl_ProductSum_for_acc_20_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_24_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_23_z);
  assign ProductSum_for_acc_20_nl = nl_ProductSum_for_acc_20_nl[34:0];
  assign nl_ProductSum_for_acc_21_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_22_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_21_z);
  assign ProductSum_for_acc_21_nl = nl_ProductSum_for_acc_21_nl[34:0];
  assign nl_ProductSum_for_acc_19_nl = ProductSum_for_acc_20_nl + ProductSum_for_acc_21_nl;
  assign ProductSum_for_acc_19_nl = nl_ProductSum_for_acc_19_nl[34:0];
  assign PECore_UpdateFSM_switch_lp_not_36_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_2_itm
      = MUX_v_35_2_2(35'b00000000000000000000000000000000000, ProductSum_for_acc_19_nl,
      PECore_UpdateFSM_switch_lp_not_36_nl);
  assign nl_ProductSum_for_acc_15_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_30_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_29_z);
  assign ProductSum_for_acc_15_nl = nl_ProductSum_for_acc_15_nl[34:0];
  assign nl_ProductSum_for_acc_13_nl = ProductSum_for_acc_14_itm_1 + ProductSum_for_acc_15_nl;
  assign ProductSum_for_acc_13_nl = nl_ProductSum_for_acc_13_nl[34:0];
  assign PECore_UpdateFSM_switch_lp_not_35_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_3_itm
      = MUX_v_35_2_2(35'b00000000000000000000000000000000000, ProductSum_for_acc_13_nl,
      PECore_UpdateFSM_switch_lp_not_35_nl);
  assign nl_ProductSum_for_acc_17_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_28_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_27_z);
  assign ProductSum_for_acc_17_nl = nl_ProductSum_for_acc_17_nl[34:0];
  assign nl_ProductSum_for_acc_18_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_26_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_25_z);
  assign ProductSum_for_acc_18_nl = nl_ProductSum_for_acc_18_nl[34:0];
  assign nl_ProductSum_for_acc_16_nl = ProductSum_for_acc_17_nl + ProductSum_for_acc_18_nl;
  assign ProductSum_for_acc_16_nl = nl_ProductSum_for_acc_16_nl[34:0];
  assign PECore_UpdateFSM_switch_lp_not_34_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_4_itm
      = MUX_v_35_2_2(35'b00000000000000000000000000000000000, ProductSum_for_acc_16_nl,
      PECore_UpdateFSM_switch_lp_not_34_nl);
  assign nl_ProductSum_for_acc_23_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_20_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_19_z);
  assign ProductSum_for_acc_23_nl = nl_ProductSum_for_acc_23_nl[34:0];
  assign nl_ProductSum_for_acc_24_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_18_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_17_z);
  assign ProductSum_for_acc_24_nl = nl_ProductSum_for_acc_24_nl[34:0];
  assign nl_ProductSum_for_acc_22_nl = ProductSum_for_acc_23_nl + ProductSum_for_acc_24_nl;
  assign ProductSum_for_acc_22_nl = nl_ProductSum_for_acc_22_nl[34:0];
  assign PECore_UpdateFSM_switch_lp_not_23_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_5_itm
      = MUX_v_35_2_2(35'b00000000000000000000000000000000000, ProductSum_for_acc_22_nl,
      PECore_UpdateFSM_switch_lp_not_23_nl);
  assign nl_ProductSum_for_acc_29_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_12_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_11_z);
  assign ProductSum_for_acc_29_nl = nl_ProductSum_for_acc_29_nl[34:0];
  assign nl_ProductSum_for_acc_30_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_10_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_9_z);
  assign ProductSum_for_acc_30_nl = nl_ProductSum_for_acc_30_nl[34:0];
  assign nl_ProductSum_for_acc_28_nl = ProductSum_for_acc_29_nl + ProductSum_for_acc_30_nl;
  assign ProductSum_for_acc_28_nl = nl_ProductSum_for_acc_28_nl[34:0];
  assign PECore_UpdateFSM_switch_lp_not_33_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_6_itm
      = MUX_v_35_2_2(35'b00000000000000000000000000000000000, ProductSum_for_acc_28_nl,
      PECore_UpdateFSM_switch_lp_not_33_nl);
  assign nl_ProductSum_for_acc_34_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_4_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_3_z);
  assign ProductSum_for_acc_34_nl = nl_ProductSum_for_acc_34_nl[34:0];
  assign nl_ProductSum_for_acc_35_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_2_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_1_z);
  assign ProductSum_for_acc_35_nl = nl_ProductSum_for_acc_35_nl[34:0];
  assign nl_ProductSum_for_acc_nl = ProductSum_for_acc_34_nl + ProductSum_for_acc_35_nl;
  assign ProductSum_for_acc_nl = nl_ProductSum_for_acc_nl[34:0];
  assign PECore_UpdateFSM_switch_lp_not_39_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_7_itm
      = MUX_v_35_2_2(35'b00000000000000000000000000000000000, ProductSum_for_acc_nl,
      PECore_UpdateFSM_switch_lp_not_39_nl);
  assign nl_ProductSum_for_acc_32_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_8_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_7_z);
  assign ProductSum_for_acc_32_nl = nl_ProductSum_for_acc_32_nl[34:0];
  assign nl_ProductSum_for_acc_33_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_6_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_5_z);
  assign ProductSum_for_acc_33_nl = nl_ProductSum_for_acc_33_nl[34:0];
  assign nl_ProductSum_for_acc_31_nl = ProductSum_for_acc_32_nl + ProductSum_for_acc_33_nl;
  assign ProductSum_for_acc_31_nl = nl_ProductSum_for_acc_31_nl[34:0];
  assign PECore_UpdateFSM_switch_lp_not_32_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_itm
      = MUX_v_35_2_2(35'b00000000000000000000000000000000000, ProductSum_for_acc_31_nl,
      PECore_UpdateFSM_switch_lp_not_32_nl);
  assign mux_59_nl = MUX_s_1_2_2(or_tmp_54, (~ mux_tmp_56), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_58_nl = MUX_s_1_2_2((~ mux_tmp_56), or_tmp_54, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_60_nl = MUX_s_1_2_2(mux_59_nl, mux_58_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_57_nl = MUX_s_1_2_2((~ mux_tmp_56), or_tmp_54, or_202_cse);
  assign mux_61_nl = MUX_s_1_2_2(mux_60_nl, mux_57_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign weight_mem_banks_load_store_for_else_and_25_ssc = PECoreRun_wen & (~ mux_61_nl)
      & and_dcpl_59;
  assign weight_port_read_out_data_and_88_enex5 = weight_port_read_out_data_and_76_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo;
  assign mux1h_4_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[15]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_15,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1[15]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[15]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[15]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[63]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63]),
      weight_port_read_out_data_0_3_sva_mx0_15, {and_929_cse , and_930_cse , and_931_cse
      , and_932_cse , and_933_cse , and_934_cse , and_935_cse , nor_397_cse});
  assign weight_port_read_out_data_0_3_sva_dfm_mx0w3_15 = mux1h_4_nl & (~ or_dcpl);
  assign mux1h_6_nl = MUX1HOT_v_15_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[14:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_14_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1[14:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[14:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[14:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[62:48]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[62:48]),
      weight_port_read_out_data_0_3_sva_mx0_14_0, {and_929_cse , and_930_cse , and_931_cse
      , and_932_cse , and_933_cse , and_934_cse , and_935_cse , nor_397_cse});
  assign not_1917_nl = ~ or_dcpl;
  assign weight_port_read_out_data_0_3_sva_dfm_mx0w3_14_0 = MUX_v_15_2_2(15'b000000000000000,
      mux1h_6_nl, not_1917_nl);
  assign weight_port_read_out_data_and_89_enex5 = weight_port_read_out_data_and_61_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_4_1_enexo;
  assign weight_mem_run_3_for_5_and_180_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_port_read_out_data_and_64_ssc = PECoreRun_wen & ((~ mux_2_itm) |
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | (~ while_stage_0_6)) & and_dcpl_48;
  assign weight_port_read_out_data_and_90_enex5 = weight_port_read_out_data_and_72_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo;
  assign and_654_ssc = and_dcpl_266 & nor_275_cse & (~ mux_259_tmp);
  assign and_656_ssc = and_dcpl_265 & while_stage_0_6 & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])
      & (~ mux_259_tmp);
  assign and_657_ssc = and_dcpl_266 & and_dcpl_643 & (~ mux_259_tmp);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_2
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 & (~ or_dcpl_316);
  assign mux1h_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[15]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1[15]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_15,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1[15]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1[15]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[15]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[15]),
      weight_port_read_out_data_0_0_sva_dfm_2_15, {crossbar_spec_PE_Weight_WordType_8U_8U_for_and_ssc
      , and_947_cse , and_948_cse , and_949_cse , and_950_cse , and_951_cse , and_952_cse
      , nor_399_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w1_15 = mux1h_nl & (~ or_dcpl_316);
  assign mux1h_9_nl = MUX1HOT_v_15_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[14:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1[14:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_14_0,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1[14:0]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1[14:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[14:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[14:0]),
      weight_port_read_out_data_0_0_sva_dfm_2_14_0, {crossbar_spec_PE_Weight_WordType_8U_8U_for_and_ssc
      , and_947_cse , and_948_cse , and_949_cse , and_950_cse , and_951_cse , and_952_cse
      , nor_399_cse});
  assign not_1921_nl = ~ or_dcpl_316;
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w1_14_0 = MUX_v_15_2_2(15'b000000000000000,
      mux1h_9_nl, not_1921_nl);
  assign weight_port_read_out_data_0_3_sva_mx0_15 = MUX1HOT_s_1_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_15,
      weight_port_read_out_data_0_3_sva_dfm_1_1_15, weight_port_read_out_data_0_3_sva_rsp_0,
      {and_dcpl_362 , and_dcpl_45 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_3_sva_mx0_14_0 = MUX1HOT_v_15_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_14_0,
      weight_port_read_out_data_0_3_sva_dfm_1_1_14_0, weight_port_read_out_data_0_3_sva_rsp_1,
      {and_dcpl_362 , and_dcpl_45 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_1_sva_mx0_15 = MUX1HOT_s_1_3_2(weight_port_read_out_data_0_1_sva_dfm_1_15,
      weight_port_read_out_data_0_1_sva_dfm_1_1_15, weight_port_read_out_data_0_1_sva_15,
      {and_dcpl_362 , and_dcpl_45 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_1_sva_mx0_14_0 = MUX1HOT_v_15_3_2(weight_port_read_out_data_0_1_sva_dfm_1_14_0,
      weight_port_read_out_data_0_1_sva_dfm_1_1_14_0, weight_port_read_out_data_0_1_sva_14_0,
      {and_dcpl_362 , and_dcpl_45 , (~ while_stage_0_8)});
  assign and_964_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_28 & (~ or_dcpl_316);
  assign mux1h_5_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1[15]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_15,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1[15]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[15]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[15]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[47]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[47]),
      weight_port_read_out_data_0_2_sva_mx0_15, {and_964_ssc , and_947_cse , and_948_cse
      , and_949_cse , and_950_cse , and_951_cse , and_952_cse , nor_399_cse});
  assign weight_port_read_out_data_0_2_sva_dfm_mx0w1_15 = mux1h_5_nl & (~ or_dcpl_316);
  assign mux1h_10_nl = MUX1HOT_v_15_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1[14:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_14_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1[14:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[14:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[14:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[46:32]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[46:32]),
      weight_port_read_out_data_0_2_sva_mx0_14_0, {and_964_ssc , and_947_cse , and_948_cse
      , and_949_cse , and_950_cse , and_951_cse , and_952_cse , nor_399_cse});
  assign not_1923_nl = ~ or_dcpl_316;
  assign weight_port_read_out_data_0_2_sva_dfm_mx0w1_14_0 = MUX_v_15_2_2(15'b000000000000000,
      mux1h_10_nl, not_1923_nl);
  assign or_12_nl = (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign mux_1_nl = MUX_s_1_2_2(or_12_nl, mux_tmp, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign weight_port_read_out_data_and_63_ssc = PECoreRun_wen & (~ mux_1_nl) & while_stage_0_7;
  assign weight_mem_run_3_for_5_and_195_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign and_1339_cse = weight_mem_run_3_for_land_1_lpi_1_dfm_3 & weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2;
  assign weight_port_read_out_data_and_91_enex5 = weight_port_read_out_data_and_74_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo;
  assign weight_port_read_out_data_and_92_enex5 = weight_port_read_out_data_and_76_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_1_1_1_enexo;
  assign weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_15 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_0_sva_dfm_2_15,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[15]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[15]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , and_1339_cse , reg_weight_mem_run_3_for_5_and_162_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_163_itm_2_cse , weight_mem_run_3_for_5_and_164_itm_2
      , reg_weight_mem_run_3_for_5_and_165_itm_2_cse , reg_weight_mem_run_3_for_5_and_166_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_167_itm_2_cse , reg_weight_mem_run_3_for_5_and_168_itm_2_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_14_0 = MUX1HOT_v_15_9_2(weight_port_read_out_data_0_0_sva_dfm_2_14_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[14:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[14:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[14:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[14:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[14:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[14:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[14:0]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[14:0]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , and_1339_cse , reg_weight_mem_run_3_for_5_and_162_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_163_itm_2_cse , weight_mem_run_3_for_5_and_164_itm_2
      , reg_weight_mem_run_3_for_5_and_165_itm_2_cse , reg_weight_mem_run_3_for_5_and_166_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_167_itm_2_cse , reg_weight_mem_run_3_for_5_and_168_itm_2_cse});
  assign weight_port_read_out_data_0_2_sva_mx0_15 = MUX1HOT_s_1_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_15,
      weight_port_read_out_data_0_2_sva_dfm_1_1_15, weight_port_read_out_data_0_2_sva_rsp_0,
      {and_dcpl_362 , and_dcpl_45 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_2_sva_mx0_14_0 = MUX1HOT_v_15_3_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0,
      weight_port_read_out_data_0_2_sva_dfm_1_1_14_0, weight_port_read_out_data_0_2_sva_rsp_1,
      {and_dcpl_362 , and_dcpl_45 , (~ while_stage_0_8)});
  assign or_tmp_320 = PECore_UpdateFSM_switch_lp_equal_tmp_2_10 | (~(PECore_RunMac_PECore_RunMac_if_and_svs_10
      | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_10)));
  assign or_688_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_2
      | reg_weight_mem_run_3_for_5_and_162_itm_2_cse | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2 | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_166_itm_2_cse | reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_2;
  assign mux_tmp_268 = MUX_s_1_2_2(or_dcpl_219, or_688_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign not_tmp_469 = ~(while_stage_0_6 | (~ mux_tmp_268));
  assign or_dcpl_325 = weight_mem_run_3_for_5_and_156_itm_2 | PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
  assign or_dcpl_336 = weight_mem_run_3_for_5_and_159_itm_2 | weight_mem_run_3_for_5_and_150_itm_2;
  assign or_dcpl_368 = weight_mem_run_3_for_5_and_95_itm_2 | weight_mem_run_3_for_5_and_86_itm_1;
  assign and_dcpl_891 = while_stage_0_3 & fsm_output;
  assign or_tmp_374 = PECore_UpdateFSM_switch_lp_equal_tmp_2_9 | (~(PECore_RunMac_PECore_RunMac_if_and_svs_9
      | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_9)));
  assign or_889_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[1])
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1;
  assign or_888_nl = (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[1]))
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1;
  assign mux_333_nl = MUX_s_1_2_2(or_889_nl, or_888_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[2]);
  assign or_887_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1;
  assign mux_334_nl = MUX_s_1_2_2(mux_333_nl, or_887_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[0]);
  assign or_tmp_406 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | mux_334_nl;
  assign or_tmp_407 = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | rva_in_reg_rw_sva_st_1_5 | (~ or_tmp_406);
  assign or_892_nl = (~ while_stage_0_8) | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1;
  assign mux_335_itm = MUX_s_1_2_2(or_892_nl, or_tmp_406, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign or_894_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_2
      | reg_weight_mem_run_3_for_5_and_162_itm_2_cse | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_166_itm_2_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2
      | reg_weight_mem_run_3_for_5_and_168_itm_2_cse;
  assign mux_tmp_323 = MUX_s_1_2_2(or_dcpl_219, or_894_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign not_tmp_653 = ~(while_stage_0_6 | (~ mux_tmp_323));
  assign nand_64_nl = ~(while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6);
  assign mux_345_nl = MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[1]),
      (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[1])), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[2]);
  assign mux_346_nl = MUX_s_1_2_2(mux_345_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse,
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[0]);
  assign or_901_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | mux_346_nl;
  assign mux_347_cse = MUX_s_1_2_2(nand_64_nl, or_901_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign not_tmp_658 = ~(while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      | mux_347_cse));
  assign or_905_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_2
      | reg_weight_mem_run_3_for_5_and_162_itm_2_cse | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_2 | reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_168_itm_2_cse;
  assign mux_tmp_335 = MUX_s_1_2_2(or_dcpl_219, or_905_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign not_tmp_662 = ~(while_stage_0_6 | (~ mux_tmp_335));
  assign or_tmp_425 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1;
  assign and_tmp_24 = while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (or_tmp_425 | mux_347_cse);
  assign data_in_tmp_operator_2_for_and_tmp = PECoreRun_wen & and_dcpl_48 & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign rva_in_reg_data_and_tmp = PECoreRun_wen & and_dcpl_292 & (and_289_cse |
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign input_mem_banks_read_1_read_data_and_4_tmp = PECoreRun_wen & (and_374_cse
      | ((~ reg_rva_in_reg_rw_sva_st_1_1_cse) & input_read_req_valid_lpi_1_dfm_1_1
      & and_dcpl_189));
  assign input_mem_banks_read_read_data_and_45_tmp = PECoreRun_wen & (~((~((~(rva_in_reg_rw_sva_st_1_4
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1))
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
      & while_stage_0_6;
  assign pe_manager_base_input_and_tmp = PECoreRun_wen & ((nand_58_cse & while_stage_0_3)
      | and_dcpl_197);
  assign and_1337_nl = weight_mem_run_3_for_land_1_lpi_1_dfm_2 & while_stage_0_6;
  assign mux_337_nl = MUX_s_1_2_2((~ mux_335_itm), or_tmp_407, and_1337_nl);
  assign and_1338_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & while_stage_0_6;
  assign mux_336_nl = MUX_s_1_2_2((~ mux_335_itm), or_tmp_407, and_1338_nl);
  assign mux_338_nl = MUX_s_1_2_2(mux_337_nl, mux_336_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_1313_tmp = (~ mux_338_nl) & and_dcpl_212 & PECoreRun_wen;
  assign accum_vector_data_and_16_cse = (~ or_dcpl_314) & fsm_output;
  assign accum_vector_data_and_17_cse = (~ or_dcpl_315) & fsm_output;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_31_cse <= 1'b0;
      reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_30_cse <= 1'b0;
      reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_7_cse <= 1'b0;
      reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_3_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_act_port_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      pe_config_manager_counter_sva_dfm_3_1 <= 4'b0000;
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= 1'b0;
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= 1'b0;
      while_stage_0_3 <= 1'b0;
      while_stage_0_4 <= 1'b0;
      while_stage_0_5 <= 1'b0;
      while_stage_0_6 <= 1'b0;
      while_stage_0_7 <= 1'b0;
      while_stage_0_8 <= 1'b0;
      while_stage_0_9 <= 1'b0;
      while_stage_0_10 <= 1'b0;
      while_stage_0_11 <= 1'b0;
      while_stage_0_12 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_164_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_145_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_133_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_5_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_4_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_1 <= 1'b0;
      input_read_addrs_sva_1_1 <= 8'b00000000;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= 1'b0;
      weight_port_read_out_data_0_3_sva_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_1_sva_15 <= 1'b0;
      weight_port_read_out_data_0_2_sva_rsp_0 <= 1'b0;
    end
    else if ( PECoreRun_wen ) begin
      reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_31_cse <= and_528_rmff;
      reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_30_cse <= and_531_rmff;
      reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_7_cse <= and_533_rmff;
      reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_3_cse <= and_534_rmff;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= and_537_rmff;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= and_539_rmff;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= and_543_rmff;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= and_546_rmff;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= and_550_rmff;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= and_554_rmff;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= and_557_rmff;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= and_560_rmff;
      reg_rva_out_Push_mioi_iswt0_cse <= and_562_cse;
      reg_start_PopNB_mioi_iswt0_cse <= and_565_rmff;
      reg_act_port_Push_mioi_iswt0_cse <= and_567_cse;
      reg_rva_in_PopNB_mioi_iswt0_cse <= fsm_output;
      pe_config_manager_counter_sva_dfm_3_1 <= MUX_v_4_2_2(4'b0000, operator_4_false_acc_nl,
          pe_config_UpdateManagerCounter_if_not_7_nl);
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= ~((pe_config_input_counter_sva_mx1 != (operator_16_false_acc_sdt_sva_1[7:0]))
          | (operator_16_false_acc_sdt_sva_1[8]));
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
      while_stage_0_3 <= reg_rva_in_PopNB_mioi_iswt0_cse;
      while_stage_0_4 <= while_stage_0_3;
      while_stage_0_5 <= while_stage_0_4;
      while_stage_0_6 <= while_stage_0_5;
      while_stage_0_7 <= while_stage_0_6;
      while_stage_0_8 <= while_stage_0_7;
      while_stage_0_9 <= while_stage_0_8;
      while_stage_0_10 <= while_stage_0_9;
      while_stage_0_11 <= while_stage_0_10;
      while_stage_0_12 <= while_stage_0_11;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_164_itm_1 <= pe_manager_base_weight_sva_mx2[2];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_145_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[1];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_133_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[0];
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1 <= ~ (pe_manager_base_weight_sva_mx2[2]);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_5_itm_1 <= ~ (pe_manager_base_weight_sva_mx1_3_0[0]);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_4_itm_1 <= ~ (pe_manager_base_weight_sva_mx1_3_0[1]);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_1
          <= ~((pe_manager_base_weight_sva_mx2[2]) | (pe_manager_base_weight_sva_mx1_3_0[1:0]!=2'b00));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1 <= (pe_manager_base_weight_sva_mx2[2])
          & (pe_manager_base_weight_sva_mx1_3_0[1:0]==2'b11) & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 <= (pe_manager_base_weight_sva_mx2[2])
          & (pe_manager_base_weight_sva_mx1_3_0[1:0]==2'b10) & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_1 <= (pe_manager_base_weight_sva_mx2[2])
          & (pe_manager_base_weight_sva_mx1_3_0[1:0]==2'b01) & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      input_read_addrs_sva_1_1 <= nl_input_read_addrs_sva_1_1[7:0];
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
      weight_port_read_out_data_0_3_sva_rsp_0 <= weight_port_read_out_data_0_3_sva_mx0_15;
      weight_port_read_out_data_0_1_sva_15 <= weight_port_read_out_data_0_1_sva_mx0_15;
      weight_port_read_out_data_0_2_sva_rsp_0 <= weight_port_read_out_data_0_2_sva_mx0_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_10 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_2_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_10 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_10 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_113_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_10 <= rva_out_reg_data_15_9_sva_dfm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_8 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_114_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_8 <= rva_out_reg_data_23_17_sva_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_8 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_115_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_8 <= rva_out_reg_data_30_25_sva_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_116_enex5 ) begin
      rva_out_reg_data_127_112_sva_dfm_4_5 <= rva_out_reg_data_127_112_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_96_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_117_enex5 ) begin
      rva_out_reg_data_111_96_sva_dfm_4_5 <= rva_out_reg_data_111_96_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_80_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_118_enex5 ) begin
      rva_out_reg_data_95_80_sva_dfm_4_5 <= rva_out_reg_data_95_80_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_119_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_4_5 <= rva_out_reg_data_79_64_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_63_sva_dfm_4_5 <= 1'b0;
      rva_out_reg_data_47_sva_dfm_4_5 <= 1'b0;
      input_read_req_valid_lpi_1_dfm_1_10 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_20_cse ) begin
      rva_out_reg_data_63_sva_dfm_4_5 <= rva_out_reg_data_63_sva_dfm_4_4;
      rva_out_reg_data_47_sva_dfm_4_5 <= rva_out_reg_data_47_sva_dfm_4_4;
      input_read_req_valid_lpi_1_dfm_1_10 <= input_read_req_valid_lpi_1_dfm_1_9;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_4_5 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_120_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_4_5 <= rva_out_reg_data_62_48_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_121_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_5 <= rva_out_reg_data_46_40_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_5 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_122_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_5 <= rva_out_reg_data_39_36_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_5 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_123_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_5 <= rva_out_reg_data_35_32_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_5_15 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_5_rsp_0 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_61_cse ) begin
      weight_port_read_out_data_0_0_sva_dfm_5_15 <= reg_weight_port_read_out_data_0_0_sva_dfm_4_ftd;
      weight_port_read_out_data_0_1_sva_dfm_5_rsp_0 <= weight_port_read_out_data_0_1_sva_dfm_4_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_5_14_0 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_78_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_5_14_0 <= reg_weight_port_read_out_data_0_0_sva_dfm_4_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_7_1_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_15_9_sva_dfm_6_6 <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_6_5_0 <= 6'b000000;
      rva_out_reg_data_23_17_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_30_25_sva_dfm_6 <= 6'b000000;
      rva_out_reg_data_0_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_8_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_16_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_31_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_24_sva_dfm_6 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_cse ) begin
      rva_out_reg_data_7_1_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_10;
      rva_out_reg_data_15_9_sva_dfm_6_6 <= PECore_PushAxiRsp_if_mux1h_12_6;
      rva_out_reg_data_15_9_sva_dfm_6_5_0 <= PECore_PushAxiRsp_if_mux1h_12_5_0;
      rva_out_reg_data_23_17_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_14;
      rva_out_reg_data_30_25_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_16;
      rva_out_reg_data_0_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_9;
      rva_out_reg_data_8_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_11;
      rva_out_reg_data_16_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_13;
      rva_out_reg_data_31_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_17;
      rva_out_reg_data_24_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_48_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_49_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_50_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_51_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_10 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
          <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_cse ) begin
      rva_in_reg_rw_sva_10 <= rva_in_reg_rw_sva_9;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_10 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_6 ) begin
      rva_in_reg_rw_sva_st_1_10 <= rva_in_reg_rw_sva_st_1_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_255_224_sva_dfm_1_1 <= 32'b00000000000000000000000000000000;
      act_port_reg_data_191_160_sva_dfm_1_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_reg_data_and_8_cse ) begin
      act_port_reg_data_255_224_sva_dfm_1_1 <= act_port_reg_data_255_224_sva_dfm_3;
      act_port_reg_data_191_160_sva_dfm_1_1 <= act_port_reg_data_191_160_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10 <= 1'b0;
      PECore_RunMac_PECore_RunMac_if_and_svs_10 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_10 <= 1'b0;
    end
    else if ( PECore_PushOutput_if_and_cse ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
      PECore_RunMac_PECore_RunMac_if_and_svs_10 <= PECore_RunMac_PECore_RunMac_if_and_svs_9;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_10 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_31_0_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_63_32_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_95_64_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_127_96_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_159_128_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_223_192_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( and_985_cse ) begin
      act_port_reg_data_31_0_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_31_0_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_27_nl);
      act_port_reg_data_63_32_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_63_32_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_28_nl);
      act_port_reg_data_95_64_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_95_64_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_29_nl);
      act_port_reg_data_127_96_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_127_96_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_30_nl);
      act_port_reg_data_159_128_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_159_128_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_31_nl);
      act_port_reg_data_223_192_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_223_192_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_19_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_10 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_28 & or_649_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_10 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_6_34_0_sva <= 35'b00000000000000000000000000000000000;
      accum_vector_data_4_34_0_sva <= 35'b00000000000000000000000000000000000;
      accum_vector_data_3_34_0_sva <= 35'b00000000000000000000000000000000000;
      accum_vector_data_2_34_0_sva <= 35'b00000000000000000000000000000000000;
      accum_vector_data_1_34_0_sva <= 35'b00000000000000000000000000000000000;
      accum_vector_data_0_34_0_sva <= 35'b00000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_8_cse ) begin
      accum_vector_data_6_34_0_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_6_itm;
      accum_vector_data_4_34_0_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_4_itm;
      accum_vector_data_3_34_0_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_3_itm;
      accum_vector_data_2_34_0_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_2_itm;
      accum_vector_data_1_34_0_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_1_itm;
      accum_vector_data_0_34_0_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_acc_14_itm_1 <= 35'b00000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_35 & PECore_RunMac_PECore_RunMac_if_and_svs_8
        & (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8) ) begin
      ProductSum_for_acc_14_itm_1 <= nl_ProductSum_for_acc_14_itm_1[34:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_35 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_8)
        ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_9 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_1_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_9 <= PECore_RunMac_PECore_RunMac_if_and_svs_8;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9
          <= 1'b0;
      rva_in_reg_rw_sva_9 <= 1'b0;
    end
    else if ( while_if_and_6_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8;
      rva_in_reg_rw_sva_9 <= rva_in_reg_rw_sva_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_34_0_sva <= 35'b00000000000000000000000000000000000;
      accum_vector_data_5_34_0_sva <= 35'b00000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_14_cse ) begin
      accum_vector_data_7_34_0_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_7_itm;
      accum_vector_data_5_34_0_sva <= PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_5_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_41 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_7)
        ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_8 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_2_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_8 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_10_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8
          <= 1'b0;
      rva_in_reg_rw_sva_8 <= 1'b0;
    end
    else if ( while_if_and_7_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_8
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
      rva_in_reg_rw_sva_8 <= rva_in_reg_rw_sva_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_45 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_6)
        ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_3_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= 1'b0;
      rva_in_reg_rw_sva_7 <= 1'b0;
      weight_port_read_out_data_0_3_sva_rsp_1 <= 15'b000000000000000;
      weight_port_read_out_data_0_1_sva_14_0 <= 15'b000000000000000;
      weight_port_read_out_data_0_2_sva_rsp_1 <= 15'b000000000000000;
    end
    else if ( while_if_and_8_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
      rva_in_reg_rw_sva_7 <= rva_in_reg_rw_sva_6;
      weight_port_read_out_data_0_3_sva_rsp_1 <= weight_port_read_out_data_0_3_sva_mx0_14_0;
      weight_port_read_out_data_0_1_sva_14_0 <= weight_port_read_out_data_0_1_sva_mx0_14_0;
      weight_port_read_out_data_0_2_sva_rsp_1 <= weight_port_read_out_data_0_2_sva_mx0_14_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_15 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_1_1_15 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_1_1_15 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_64_ssc ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_15 <= MUX1HOT_s_1_9_2(weight_port_read_out_data_0_2_sva_mx0_15,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[31]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55
          , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_185_ssc , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_179_cse , weight_mem_run_3_for_5_and_188_cse
          , weight_mem_run_3_for_5_and_189_ssc});
      weight_port_read_out_data_0_1_sva_dfm_1_1_15 <= MUX1HOT_s_1_9_2(weight_port_read_out_data_0_1_sva_mx0_15,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[31]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[15]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55
          , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_179_cse , weight_mem_run_3_for_5_and_180_ssc
          , weight_mem_run_3_for_5_and_181_cse});
      weight_port_read_out_data_0_3_sva_dfm_1_1_15 <= MUX1HOT_s_1_9_2(weight_port_read_out_data_0_3_sva_mx0_15,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[47]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55
          , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_195_ssc , weight_mem_run_3_for_5_and_188_cse
          , weight_mem_run_3_for_5_and_181_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_14_0 <= 15'b000000000000000;
    end
    else if ( mux_287_nl & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & while_stage_0_7 & PECoreRun_wen ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1_14_0 <= MUX1HOT_v_15_9_2(weight_port_read_out_data_0_2_sva_mx0_14_0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[46:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[46:32]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[46:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[46:32]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[46:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[46:32]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[46:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[30:16]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55
          , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_185_ssc , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_179_cse , weight_mem_run_3_for_5_and_188_cse
          , weight_mem_run_3_for_5_and_189_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_5_mux_4_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_5_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_6_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_7_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_48_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_49_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_50_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_51_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_52_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_53_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_54_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_55_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_8_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_9_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_14_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_23_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_32_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_33_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_34_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_35_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_36_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_37_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_38_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_39_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_24_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_25_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_26_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_27_itm_1 <= 16'b0000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_cse ) begin
      weight_mem_run_3_for_5_mux_4_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_4_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_5_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_5_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_6_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_6_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_7_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_7_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_48_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_49_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_1_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_50_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_51_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_52_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_53_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_54_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_55_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_8_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_9_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_1_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_14_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000006,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_23_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_2_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_3_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_32_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_4_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_33_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_4_1_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_34_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_4_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_35_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_4_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_36_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_4_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_37_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_4_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_38_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_4_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_39_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_4_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_24_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_25_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_1_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_26_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_27_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_7_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_enex5 ) begin
      weight_port_read_out_data_1_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
          <= 16'b0000000000000000;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
          <= MUX_v_16_2_2(16'b0000000000000000, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_2_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= 1'b0;
      rva_in_reg_rw_sva_6 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_cse ) begin
      weight_mem_run_3_for_land_2_lpi_1_dfm_3 <= weight_mem_run_3_for_land_2_lpi_1_dfm_2;
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= weight_mem_run_3_for_land_3_lpi_1_dfm_2;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
      rva_in_reg_rw_sva_6 <= rva_in_reg_rw_sva_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_79_enex5 ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000005
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000004
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000006
          <= 16'b0000000000000000;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[15:0]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[31:16]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[47:32]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000005
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[63:48]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000004
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[79:64]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000006
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[95:80]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_80_enex5 ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_81_enex5 ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_3_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_82_enex5 ) begin
      weight_port_read_out_data_2_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_4_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_83_enex5 ) begin
      weight_port_read_out_data_2_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000005;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_5_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_84_enex5 ) begin
      weight_port_read_out_data_2_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000004;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_6_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_85_enex5 ) begin
      weight_port_read_out_data_2_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_4_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_5,
          weight_port_read_out_data_0_3_sva_dfm_mx0w3_15, PECore_PushAxiRsp_if_else_mux_18_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_30_tmp , while_and_29_cse});
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5,
          weight_port_read_out_data_0_2_sva_dfm_mx0w1_15, PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_30_tmp , while_and_29_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        & while_stage_0_6 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        & while_stage_0_6 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_5 <= 1'b0;
      weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6 <= 2'b00;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3 <= 3'b000;
      rva_in_reg_rw_sva_st_5 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_2_cse ) begin
      rva_in_reg_rw_sva_st_1_5 <= rva_in_reg_rw_sva_st_1_4;
      weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6 <= weight_mem_write_arbxbar_xbar_for_empty_sva_2[7:6];
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
      rva_in_reg_rw_sva_st_5 <= rva_in_reg_rw_sva_st_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_1_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_2 <= 1'b0;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= 1'b0;
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_run_3_for_5_and_156_itm_2 <= 1'b0;
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_run_3_for_5_and_159_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_2 <= 1'b0;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2 <= 1'b0;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_92_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_94_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_95_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_86_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_88_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_71_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_7_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_60_itm_1 <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_30_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_31_itm_1 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_20_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_15_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_8_itm_1 <= 1'b0;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_162_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_163_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_164_itm_2 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_165_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_166_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_167_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_168_itm_2_cse <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_5_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_run_3_for_5_and_156_itm_2 <= weight_mem_run_3_for_5_and_156_itm_1;
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= MUX_v_128_2_2(weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_run_3_for_5_and_159_itm_2 <= weight_mem_run_3_for_5_and_159_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_2_2_0!=3'b000));
      weight_mem_run_3_for_5_and_150_itm_2 <= weight_mem_run_3_for_5_and_150_itm_1;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= weight_read_addrs_7_lpi_1_dfm_2_2_0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_1;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_92_itm_2 <= weight_mem_run_3_for_5_and_92_itm_1;
      weight_mem_run_3_for_5_and_94_itm_2 <= weight_mem_run_3_for_5_and_94_itm_1;
      weight_mem_run_3_for_5_and_95_itm_2 <= weight_mem_run_3_for_5_and_95_itm_1;
      weight_mem_run_3_for_5_and_86_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b101)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_88_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b111)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_71_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b110)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_7_itm_1 <= ~((weight_read_addrs_5_lpi_1_dfm_2_2_0!=3'b000));
      weight_mem_run_3_for_5_and_60_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b011)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= weight_read_addrs_5_lpi_1_dfm_2_2_0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1_1;
      reg_weight_mem_run_3_for_5_and_30_itm_2_cse <= weight_mem_run_3_for_5_and_30_itm_1;
      weight_mem_run_3_for_5_and_31_itm_1 <= (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b110)
          & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
      reg_weight_mem_run_3_for_5_and_20_itm_2_cse <= weight_mem_run_3_for_5_and_20_itm_1;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
      reg_weight_mem_run_3_for_5_and_15_itm_2_cse <= weight_mem_run_3_for_5_and_15_itm_1;
      weight_mem_run_3_for_5_and_8_itm_1 <= (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b111)
          & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= weight_read_addrs_3_lpi_1_dfm_2_2_0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1;
      reg_weight_mem_run_3_for_5_and_162_itm_2_cse <= weight_mem_run_3_for_5_and_162_itm_1;
      reg_weight_mem_run_3_for_5_and_163_itm_2_cse <= weight_mem_run_3_for_5_and_163_itm_1;
      weight_mem_run_3_for_5_and_164_itm_2 <= weight_mem_run_3_for_5_and_164_itm_1;
      reg_weight_mem_run_3_for_5_and_165_itm_2_cse <= weight_mem_run_3_for_5_and_165_itm_1;
      reg_weight_mem_run_3_for_5_and_166_itm_2_cse <= weight_mem_run_3_for_5_and_166_itm_1;
      reg_weight_mem_run_3_for_5_and_167_itm_2_cse <= weight_mem_run_3_for_5_and_167_itm_1;
      reg_weight_mem_run_3_for_5_and_168_itm_2_cse <= weight_mem_run_3_for_5_and_168_itm_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_7_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1053_cse | weight_mem_run_3_for_5_and_159_itm_2 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5
        | or_dcpl_325) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & while_stage_0_7 & PECoreRun_wen ) begin
      weight_port_read_out_data_7_7_sva_dfm_1 <= weight_port_read_out_data_7_7_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_6_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (((mux_289_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1)
        & weight_mem_run_3_for_land_lpi_1_dfm_2) | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5
        | weight_mem_run_3_for_5_and_150_itm_2 | or_dcpl_325) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & while_stage_0_7 & PECoreRun_wen ) begin
      weight_port_read_out_data_7_6_sva_dfm_1 <= weight_port_read_out_data_7_6_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_5_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_7_3_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_7_2_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_7_1_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( and_1062_cse ) begin
      weight_port_read_out_data_7_5_sva_dfm_1 <= weight_port_read_out_data_7_5_sva_dfm_2;
      weight_port_read_out_data_7_3_sva_dfm_1 <= weight_port_read_out_data_7_3_sva_dfm_2;
      weight_port_read_out_data_7_2_sva_dfm_1 <= weight_port_read_out_data_7_2_sva_dfm_2;
      weight_port_read_out_data_7_1_sva_dfm_1 <= weight_port_read_out_data_7_1_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_4_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_7_0_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( and_1066_cse ) begin
      weight_port_read_out_data_7_4_sva_dfm_1 <= weight_port_read_out_data_7_4_sva_dfm_2;
      weight_port_read_out_data_7_0_sva_dfm_1 <= weight_port_read_out_data_7_0_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_7_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_2_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( and_1086_cse ) begin
      weight_port_read_out_data_5_7_sva_dfm_1 <= weight_port_read_out_data_5_7_sva_dfm_2;
      weight_port_read_out_data_5_2_sva_dfm_1 <= weight_port_read_out_data_5_2_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_6_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_5_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_1_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( and_1090_cse ) begin
      weight_port_read_out_data_5_6_sva_dfm_1 <= weight_port_read_out_data_5_6_sva_dfm_2;
      weight_port_read_out_data_5_5_sva_dfm_1 <= weight_port_read_out_data_5_5_sva_dfm_2;
      weight_port_read_out_data_5_1_sva_dfm_1 <= weight_port_read_out_data_5_1_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_4_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1085_cse | weight_mem_run_3_for_5_and_71_itm_1 | weight_mem_run_3_for_5_and_86_itm_1
        | weight_mem_run_3_for_5_and_92_itm_2) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & while_stage_0_7 & PECoreRun_wen ) begin
      weight_port_read_out_data_5_4_sva_dfm_1 <= weight_port_read_out_data_5_4_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_3_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (((xor_5_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_7_itm_1)
        & weight_mem_run_3_for_land_6_lpi_1_dfm_2) | or_dcpl_368 | weight_mem_run_3_for_5_and_60_itm_1)
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & while_stage_0_7 & PECoreRun_wen ) begin
      weight_port_read_out_data_5_3_sva_dfm_1 <= weight_port_read_out_data_5_3_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (((mux_307_nl | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_7_itm_1)
        & weight_mem_run_3_for_land_6_lpi_1_dfm_2) | or_dcpl_368) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & while_stage_0_7 & PECoreRun_wen ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= weight_port_read_out_data_5_0_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_28_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_22_itm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= 1'b0;
      rva_in_reg_rw_sva_5 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_4_cse ) begin
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_28_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      weight_mem_run_3_for_5_and_22_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= weight_mem_run_3_for_land_1_lpi_1_dfm_2;
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= weight_mem_run_3_for_land_7_lpi_1_dfm_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= weight_mem_run_3_for_land_3_lpi_1_dfm_1;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= weight_mem_run_3_for_land_5_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
      rva_in_reg_rw_sva_5 <= rva_in_reg_rw_sva_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_7_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1118_cse | weight_mem_run_3_for_5_and_31_itm_1 | reg_weight_mem_run_3_for_5_and_30_itm_2_cse
        | weight_mem_run_3_for_5_and_28_itm_1) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_3_7_sva_dfm_1 <= weight_port_read_out_data_3_7_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_6_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1118_cse | weight_mem_run_3_for_5_and_31_itm_1 | weight_mem_run_3_for_5_and_22_itm_1
        | reg_weight_mem_run_3_for_5_and_20_itm_2_cse) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_3_6_sva_dfm_1 <= weight_port_read_out_data_3_6_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_5_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (((xor_13_cse | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse)
        & weight_mem_run_3_for_land_4_lpi_1_dfm_2) | reg_weight_mem_run_3_for_5_and_15_itm_2_cse
        | reg_weight_mem_run_3_for_5_and_30_itm_2_cse | reg_weight_mem_run_3_for_5_and_20_itm_2_cse)
        & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_3_5_sva_dfm_1 <= weight_port_read_out_data_3_5_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_4_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (((mux_309_nl | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse)
        & weight_mem_run_3_for_land_4_lpi_1_dfm_2) | weight_mem_run_3_for_5_and_8_itm_1
        | weight_mem_run_3_for_5_and_31_itm_1 | reg_weight_mem_run_3_for_5_and_30_itm_2_cse
        | reg_weight_mem_run_3_for_5_and_20_itm_2_cse) & fsm_output & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_3_4_sva_dfm_1 <= weight_port_read_out_data_3_4_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= 16'b0000000000000000;
    end
    else if ( (weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & while_stage_0_7 & PECoreRun_wen ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & mux_4_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1
          <= MUX_v_16_2_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[15:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & mux_5_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_128U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1
          <= MUX_v_16_2_2((weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[15:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_16 <= 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_222 | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & mux_6_nl ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_127_16 <= weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_222 | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & mux_9_nl ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_RunFSM_switch_lp_equal_tmp_1_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_UpdateFSM_switch_lp_equal_tmp_2_3 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_empty_sva_1[2])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_10_nl) & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_71 & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1 <= 1'b0;
    end
    else if ( weight_read_addrs_and_3_cse ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_22_itm_1 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_71 & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_71 & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= 1'b0;
      rva_in_reg_rw_sva_4 <= 1'b0;
    end
    else if ( while_if_and_11_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= weight_mem_run_3_for_weight_mem_run_3_for_and_3_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & or_260_cse;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & weight_mem_read_arbxbar_xbar_1_for_3_8_for_5_or_cse;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & or_253_cse;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
      rva_in_reg_rw_sva_4 <= rva_in_reg_rw_sva_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_53_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_59_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_65_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_71_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_77_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_83_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_89_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva <= 15'b000000000000000;
    end
    else if ( (~ mux_311_nl) & fsm_output & while_stage_0_5 & PECoreRun_wen ) begin
      pe_manager_base_weight_sva <= pe_manager_base_weight_sva_mx2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= 11'b00000000000;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= 1'b0;
    end
    else if ( weight_read_addrs_and_5_cse ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= MUX_v_11_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl,
          weight_read_addrs_0_14_4_lpi_1_dfm_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= MUX_s_1_2_2((weight_read_addrs_0_3_0_lpi_1_dfm_4[3]),
          (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_146 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_146 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_24_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_25_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_26_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_27_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_28_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_29_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_30_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_31_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= 12'b000000000000;
    end
    else if ( weight_write_addrs_and_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= weight_write_addrs_lpi_1_dfm_1_2[14:3];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1,
          Arbiter_8U_Roundrobin_pick_1_if_1_and_5_tmp, Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1,
          Arbiter_8U_Roundrobin_pick_1_if_1_and_8_tmp, Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_1_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_3_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= 13'b0000000000000;
      weight_read_addrs_5_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_7_lpi_1_dfm_1 <= 15'b000000000000000;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= 1'b0;
    end
    else if ( weight_read_addrs_and_7_cse ) begin
      weight_read_addrs_1_lpi_1_dfm_1 <= weight_read_addrs_1_lpi_1_dfm_1_1;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_3_lpi_1_dfm_1 <= weight_read_addrs_3_lpi_1_dfm_1_1;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_1 <= weight_read_addrs_5_lpi_1_dfm_1_1;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_7_lpi_1_dfm_1 <= weight_read_addrs_7_lpi_1_dfm_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_5_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_8_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_not_185,
          weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0, and_dcpl_580);
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0, and_108_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0, and_115_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0, and_122_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0,
          (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp);
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0, and_129_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0, and_dcpl_618);
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0,
          (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1 <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= 1'b0;
      rva_in_reg_rw_sva_3 <= 1'b0;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1 <= MUX_s_1_2_2((pe_manager_base_weight_sva_mx1_3_0[1]),
          reg_rva_in_reg_rw_sva_2_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      rva_in_reg_rw_sva_3 <= reg_rva_in_reg_rw_sva_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_31_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= 1'b0;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= 8'b00000000;
      rva_in_reg_rw_sva_st_3 <= 1'b0;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_1_for_and_cse ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_31_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b101)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b110)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= weight_mem_write_arbxbar_xbar_for_lshift_tmp;
      rva_in_reg_rw_sva_st_3 <= reg_rva_in_reg_rw_sva_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_and_cse ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_582);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_582);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_582);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_582);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_582);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_582);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_582);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_582);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_64_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse & ((~ while_stage_0_5) | while_and_1145_itm_1)
        ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= MUX_v_15_2_2(pe_manager_base_weight_sva_mx2,
          PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1, while_and_1145_itm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_32_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_7_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_33_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_6_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_34_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_5_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_35_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_36_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_3_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_37_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_2_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_38_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_1_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_39_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= 15'b000000000000000;
    end
    else if ( weight_write_addrs_and_3_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= weight_write_addrs_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( weight_write_data_data_and_8_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_2_cse <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= 1'b0;
      while_and_1145_itm_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_3_cse ) begin
      reg_rva_in_reg_rw_sva_2_cse <= reg_rva_in_reg_rw_sva_st_1_1_cse;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= MUX_s_1_2_2(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
      while_and_1145_itm_1 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1
          & PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
          & reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= 4'b0000;
    end
    else if ( weight_read_addrs_and_29_enex5 ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= 11'b00000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_193 ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_2_1_sva <= 2'b00;
      pe_config_is_zero_first_sva <= 1'b0;
    end
    else if ( state_and_cse ) begin
      state_2_1_sva <= state_mux_1_cse;
      pe_config_is_zero_first_sva <= pe_config_is_zero_first_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_0_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_226) ) begin
      state_0_sva <= PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_manager_counter_sva <= 4'b0000;
    end
    else if ( mux_312_nl & rva_in_reg_rw_and_3_cse ) begin
      pe_config_manager_counter_sva <= pe_config_manager_counter_sva_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_num_manager_sva <= 4'b0001;
      pe_config_num_output_sva <= 8'b00000001;
    end
    else if ( pe_config_num_manager_and_cse ) begin
      pe_config_num_manager_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[35:32];
      pe_config_num_output_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= 1'b0;
      state_2_1_sva_dfm_1 <= 2'b00;
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= 8'b00000000;
      input_write_req_valid_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_4_cse ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= rva_in_PopNB_mioi_return_rsc_z_mxwt;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
      state_2_1_sva_dfm_1 <= MUX_v_2_2_2(PECore_UpdateFSM_switch_lp_and_1_nl, state_mux_1_cse,
          rva_in_PopNB_mioi_return_rsc_z_mxwt);
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= and_289_cse;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0];
      input_write_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= 1'b0;
      PECore_RunFSM_switch_lp_nor_tmp_1 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_11_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= PECore_UpdateFSM_switch_lp_equal_tmp_6;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= ~(PECore_RunScale_PECore_RunScale_if_and_1_svs_1
          | PECore_UpdateFSM_switch_lp_nor_tmp_1);
      PECore_RunFSM_switch_lp_nor_tmp_1 <= ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
          | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(or_tmp_129 | or_dcpl_226)) ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= input_port_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva <= 8'b00000000;
    end
    else if ( or_804_cse & mux_313_nl & and_dcpl_891 & PECoreRun_wen ) begin
      pe_config_input_counter_sva <= pe_config_input_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva <= 8'b00000000;
    end
    else if ( or_804_cse & mux_314_nl & and_dcpl_891 & PECoreRun_wen ) begin
      pe_config_output_counter_sva <= pe_config_output_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      operator_8_false_acc_sdt_sva_1 <= 9'b000000000;
    end
    else if ( pe_config_UpdateManagerCounter_if_if_and_enex5 ) begin
      operator_8_false_acc_sdt_sva_1 <= nl_operator_8_false_acc_sdt_sva_1[8:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_manager_counter_sva_dfm_1 <= 4'b0000;
      pe_config_output_counter_sva_dfm_1 <= 8'b00000000;
      pe_config_input_counter_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1173_cse ) begin
      pe_config_manager_counter_sva_dfm_1 <= MUX_v_4_2_2(4'b0000, pe_config_manager_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
      pe_config_output_counter_sva_dfm_1 <= MUX_v_8_2_2(8'b00000000, pe_config_output_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
      pe_config_input_counter_sva_dfm_1 <= MUX_v_8_2_2(8'b00000000, pe_config_input_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiWrite_switch_lp_and_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_191_160_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_255_224_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( and_1179_cse ) begin
      act_port_reg_data_191_160_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_191_160_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_38_nl);
      act_port_reg_data_255_224_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_255_224_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_21_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & and_dcpl_216 ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & (and_dcpl_216 | and_dcpl_220) ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2 <= 2'b00;
    end
    else if ( weight_read_addrs_and_16_cse ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2 <= pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & and_dcpl_220 ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_4_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_5_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_6_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_7_sva_dfm_2 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_28_cse ) begin
      weight_port_read_out_data_0_4_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_63_48_sva_1,
          while_and_30_tmp);
      weight_port_read_out_data_0_5_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_79_64_sva_1,
          while_and_30_tmp);
      weight_port_read_out_data_0_6_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_95_80_sva_1,
          while_and_30_tmp);
      weight_port_read_out_data_0_7_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_128_127_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_16_15_0_sdt_111_96_sva_1,
          while_and_30_tmp);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_1_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_32_cse ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_6_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_1_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_2_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_3_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_4_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_5_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_6_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_40_cse ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_1_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001;
      weight_port_read_out_data_1_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002;
      weight_port_read_out_data_1_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003;
      weight_port_read_out_data_1_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000004;
      weight_port_read_out_data_1_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000005;
      weight_port_read_out_data_1_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_7_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_222 | (~ weight_mem_run_3_for_land_3_lpi_1_dfm_2)))
        ) begin
      weight_port_read_out_data_2_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_4_1_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_4_2_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_4_3_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_4_4_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_4_5_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_4_6_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_4_7_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_48_cse ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_4_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_4_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_4_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_4_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_4_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_4_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_4_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_0_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_1_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_2_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_3_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_68_cse ) begin
      weight_port_read_out_data_3_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000000;
      weight_port_read_out_data_3_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000001;
      weight_port_read_out_data_3_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002;
      weight_port_read_out_data_3_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_2
          <= MUX_s_1_2_2(weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_35_nl & while_stage_0_6 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_103_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_108_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_2_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_20_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_24_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_2 <= 1'b0;
      weight_read_addrs_1_lpi_1_dfm_3_2_0 <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_109_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_1;
      weight_read_addrs_1_lpi_1_dfm_3_2_0 <= weight_read_addrs_1_lpi_1_dfm_2_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_3
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_3 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_3 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_3 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_3
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= 1'b0;
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_5_and_159_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_156_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_95_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_94_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_92_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_30_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_20_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_15_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_168_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_167_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_166_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_165_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_164_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_163_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_162_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= 1'b0;
    end
    else if ( weight_read_addrs_and_19_cse ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= weight_read_addrs_7_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= weight_read_addrs_5_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= weight_read_addrs_3_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_5_and_159_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_156_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_150_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_95_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b110)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_94_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b101)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_92_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_1 <= ~((weight_read_addrs_5_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_30_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1;
      weight_mem_run_3_for_5_and_20_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1;
      weight_mem_run_3_for_5_and_15_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= ~((weight_read_addrs_3_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_168_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1_1;
      weight_mem_run_3_for_5_and_167_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b110)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_166_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1_1;
      weight_mem_run_3_for_5_and_165_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
      weight_mem_run_3_for_5_and_164_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1
          & (pe_manager_base_weight_sva[0]) & (~ (pe_manager_base_weight_sva[2]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_163_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
      weight_mem_run_3_for_5_and_162_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1 <= ~((pe_manager_base_weight_sva[2])
          | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1 | (pe_manager_base_weight_sva[0]));
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_36_nl ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_37_nl ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_38_nl ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        | (~ while_stage_0_6))) ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & ((~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_55_nl ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_24_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_30_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= 1'b0;
    end
    else if ( operator_15_false_1_and_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        | (~ while_stage_0_4))) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_dcpl_618 | or_dcpl_60)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_129_cse | or_dcpl_60)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        | (~ while_stage_0_4))) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_122_cse | or_dcpl_60)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_115_cse | or_dcpl_60)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_108_cse | or_dcpl_60)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= 15'b000000000000000;
    end
    else if ( PEManager_15U_PEManagerWrite_and_enex5 ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= rva_in_reg_data_sva_1[30:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_num_input_sva <= 8'b00000001;
      pe_manager_base_bias_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_num_input_and_cse ) begin
      pe_manager_num_input_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      pe_manager_base_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[46:32];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_is_valid_sva <= 1'b0;
      pe_config_is_cluster_sva <= 1'b0;
      pe_config_is_bias_sva <= 1'b0;
    end
    else if ( pe_config_is_valid_and_cse ) begin
      pe_config_is_valid_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
      pe_config_is_cluster_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[16];
      pe_config_is_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_zero_active_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & and_289_cse & (~ PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)
        & (~ or_dcpl_231) ) begin
      pe_manager_zero_active_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_mux_19_itm_1 <= 1'b0;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= 4'b0000;
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_addrs_lpi_1_dfm_1_1 <= 15'b000000000000000;
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= 11'b00000000000;
    end
    else if ( while_if_and_15_cse ) begin
      while_if_mux_19_itm_1 <= MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_19_nl,
          rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:0])
          & ({{3{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_4_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:112])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:96])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:80])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:64])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:48])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:32])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:16])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:0])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_addrs_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:0])
          & ({{14{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{14{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:4])
          & ({{10{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_11_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_48 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_5)
        ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_4 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= 3'b000;
      rva_in_reg_rw_sva_st_4 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_5_cse ) begin
      rva_in_reg_rw_sva_st_1_4 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1;
      rva_in_reg_rw_sva_st_4 <= rva_in_reg_rw_sva_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_9 <= 1'b0;
      rva_in_reg_rw_sva_st_9 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_6_cse ) begin
      rva_in_reg_rw_sva_st_1_9 <= rva_in_reg_rw_sva_st_1_8;
      rva_in_reg_rw_sva_st_9 <= rva_in_reg_rw_sva_st_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= 4'b0000;
    end
    else if ( PECoreRun_wen & and_dcpl_238 ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_9_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_52_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_53_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_54_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_55_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_17_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_2_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_9 <= 1'b0;
      rva_out_reg_data_47_sva_dfm_4_4 <= 1'b0;
      rva_out_reg_data_63_sva_dfm_4_4 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( input_read_req_valid_and_1_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_9 <= input_read_req_valid_lpi_1_dfm_1_8;
      rva_out_reg_data_47_sva_dfm_4_4 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      rva_out_reg_data_63_sva_dfm_4_4 <= PECore_RunMac_PECore_RunMac_if_and_svs_8;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_7_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_124_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= rva_out_reg_data_30_25_sva_dfm_6_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_7 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_125_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_7 <= rva_out_reg_data_23_17_sva_dfm_6_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_126_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= rva_out_reg_data_15_9_sva_dfm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_4_ftd <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_4_15 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_72_cse ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_4_ftd <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
      weight_port_read_out_data_0_1_sva_dfm_4_15 <= reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_4_ftd_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_86_enex5 ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_4_ftd_1 <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_127_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= rva_out_reg_data_35_32_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_128_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_4 <= rva_out_reg_data_39_36_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_129_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_4 <= rva_out_reg_data_46_40_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_4_4 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_130_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_4_4 <= rva_out_reg_data_62_48_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_131_enex5 ) begin
      rva_out_reg_data_127_112_sva_dfm_4_4 <= rva_out_reg_data_127_112_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_96_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_132_enex5 ) begin
      rva_out_reg_data_111_96_sva_dfm_4_4 <= rva_out_reg_data_111_96_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_80_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_133_enex5 ) begin
      rva_out_reg_data_95_80_sva_dfm_4_4 <= rva_out_reg_data_95_80_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_134_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_4_4 <= rva_out_reg_data_79_64_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_39_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_37_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_36_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= 16'b0000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_129_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_101_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_115_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_122_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_39_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_94_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_108_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_130_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_102_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_116_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_123_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_95_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_109_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_131_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_103_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_117_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_124_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_37_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_96_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_110_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_132_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_104_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_118_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_125_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_36_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_97_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_111_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1
          <= 16'b0000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_24_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[63:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_133_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[47:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & mux_63_nl & and_dcpl_266 ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, mux1h_2_nl, not_1864_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= 16'b0000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_27_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[63:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_126_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[47:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_127_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[31:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_128_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= 16'b0000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_28_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[63:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_112_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[31:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_114_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & (~ mux_81_nl) & while_stage_0_6 ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, mux_275_nl, nor_398_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_1
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        & while_stage_0_6 ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[47:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_113_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_266 & crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse
        ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[15:0]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_78_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_1_lpi_1_dfm_2_2_0 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1
          <= 1'b0;
    end
    else if ( weight_read_addrs_and_24_cse ) begin
      weight_read_addrs_1_lpi_1_dfm_2_2_0 <= weight_read_addrs_1_lpi_1_dfm_1[2:0];
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1
          <= ~((weight_read_addrs_1_lpi_1_dfm_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_data_sva_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rva_in_reg_data_and_tmp ) begin
      rva_in_reg_data_sva_1 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
        & while_stage_0_6 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]))) & while_stage_0_4 )
        begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_8 <= 1'b0;
      rva_in_reg_rw_sva_st_8 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_9_cse ) begin
      rva_in_reg_rw_sva_st_1_8 <= rva_in_reg_rw_sva_st_1_7;
      rva_in_reg_rw_sva_st_8 <= rva_in_reg_rw_sva_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse
        | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1)
        | (or_dcpl_28 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1) | (or_dcpl_42
        & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1) | ((Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1
        | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1)
        | (or_dcpl_35 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1) | (or_dcpl_53
        & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1) | ((Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1
        | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1)
        | ((Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5)
        & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)) & and_dcpl_279 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_1 <= pe_manager_base_weight_sva[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_1 <= 2'b00;
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= 1'b0;
    end
    else if ( pe_manager_base_weight_and_5_cse ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_1 <= pe_manager_base_weight_sva[1:0];
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= weight_read_addrs_4_14_2_lpi_1_dfm_1[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_117_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_31_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_122_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_38_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_83_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_164_itm_1
          & (pe_manager_base_weight_sva[1:0]==2'b10) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b011)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_6_itm_1
          <= ~((pe_manager_base_weight_sva[2:0]!=3'b000));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_1 <= (pe_manager_base_weight_sva[2])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_145_itm_1 & (pe_manager_base_weight_sva[0])
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_1 <= (pe_manager_base_weight_sva[1])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_133_itm_1 & (~
          (pe_manager_base_weight_sva[2])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_164_itm_1
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_133_itm_1 & (~
          (pe_manager_base_weight_sva[1])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_145_itm_1
          & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_89_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_nl,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1_1,
          PECore_UpdateFSM_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_nl,
          PECore_RunFSM_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_85_nl & while_stage_0_5 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_nl,
          input_read_req_valid_lpi_1_dfm_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_18_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_56_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_57_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_58_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_59_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_18_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & or_253_cse & and_dcpl_279 ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & or_260_cse & and_dcpl_279 ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( input_read_req_valid_and_2_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= input_read_req_valid_lpi_1_dfm_1_7;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_11_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_6_1 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_135_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_6_1 <= rva_out_reg_data_30_25_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_6_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_136_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_6_1 <= rva_out_reg_data_23_17_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_137_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= rva_out_reg_data_15_9_sva_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_74_cse ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd <= weight_port_read_out_data_0_1_sva_dfm_2_rsp_0;
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_0_sva_dfm_2_15_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_87_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1 <= weight_port_read_out_data_0_1_sva_dfm_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_138_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= rva_out_reg_data_35_32_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_139_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_3 <= rva_out_reg_data_39_36_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_140_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3 <= rva_out_reg_data_46_40_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_4_3 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_141_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_4_3 <= rva_out_reg_data_62_48_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_142_enex5 ) begin
      rva_out_reg_data_127_112_sva_dfm_4_3 <= rva_out_reg_data_127_112_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_96_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_143_enex5 ) begin
      rva_out_reg_data_111_96_sva_dfm_4_3 <= rva_out_reg_data_111_96_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_80_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_144_enex5 ) begin
      rva_out_reg_data_95_80_sva_dfm_4_3 <= rva_out_reg_data_95_80_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_145_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_4_3 <= rva_out_reg_data_79_64_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= 8'b00000000;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_empty_and_enex5 ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= weight_mem_write_arbxbar_xbar_for_empty_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_7_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_7 <= 1'b0;
      rva_in_reg_rw_sva_st_7 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_12_cse ) begin
      rva_in_reg_rw_sva_st_1_7 <= rva_in_reg_rw_sva_st_1_6;
      rva_in_reg_rw_sva_st_7 <= rva_in_reg_rw_sva_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_27_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_60_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_61_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_62_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_63_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= MUX_v_128_256_2(input_mem_banks_bank_a_0_sva_dfm_2,
          input_mem_banks_bank_a_1_sva_dfm_2, input_mem_banks_bank_a_2_sva_dfm_2,
          input_mem_banks_bank_a_3_sva_dfm_2, input_mem_banks_bank_a_4_sva_dfm_2,
          input_mem_banks_bank_a_5_sva_dfm_2, input_mem_banks_bank_a_6_sva_dfm_2,
          input_mem_banks_bank_a_7_sva_dfm_2, input_mem_banks_bank_a_8_sva_dfm_2,
          input_mem_banks_bank_a_9_sva_dfm_2, input_mem_banks_bank_a_10_sva_dfm_2,
          input_mem_banks_bank_a_11_sva_dfm_2, input_mem_banks_bank_a_12_sva_dfm_2,
          input_mem_banks_bank_a_13_sva_dfm_2, input_mem_banks_bank_a_14_sva_dfm_2,
          input_mem_banks_bank_a_15_sva_dfm_2, input_mem_banks_bank_a_16_sva_dfm_2,
          input_mem_banks_bank_a_17_sva_dfm_2, input_mem_banks_bank_a_18_sva_dfm_2,
          input_mem_banks_bank_a_19_sva_dfm_2, input_mem_banks_bank_a_20_sva_dfm_2,
          input_mem_banks_bank_a_21_sva_dfm_2, input_mem_banks_bank_a_22_sva_dfm_2,
          input_mem_banks_bank_a_23_sva_dfm_2, input_mem_banks_bank_a_24_sva_dfm_2,
          input_mem_banks_bank_a_25_sva_dfm_2, input_mem_banks_bank_a_26_sva_dfm_2,
          input_mem_banks_bank_a_27_sva_dfm_2, input_mem_banks_bank_a_28_sva_dfm_2,
          input_mem_banks_bank_a_29_sva_dfm_2, input_mem_banks_bank_a_30_sva_dfm_2,
          input_mem_banks_bank_a_31_sva_dfm_2, input_mem_banks_bank_a_32_sva_dfm_2,
          input_mem_banks_bank_a_33_sva_dfm_2, input_mem_banks_bank_a_34_sva_dfm_2,
          input_mem_banks_bank_a_35_sva_dfm_2, input_mem_banks_bank_a_36_sva_dfm_2,
          input_mem_banks_bank_a_37_sva_dfm_2, input_mem_banks_bank_a_38_sva_dfm_2,
          input_mem_banks_bank_a_39_sva_dfm_2, input_mem_banks_bank_a_40_sva_dfm_2,
          input_mem_banks_bank_a_41_sva_dfm_2, input_mem_banks_bank_a_42_sva_dfm_2,
          input_mem_banks_bank_a_43_sva_dfm_2, input_mem_banks_bank_a_44_sva_dfm_2,
          input_mem_banks_bank_a_45_sva_dfm_2, input_mem_banks_bank_a_46_sva_dfm_2,
          input_mem_banks_bank_a_47_sva_dfm_2, input_mem_banks_bank_a_48_sva_dfm_2,
          input_mem_banks_bank_a_49_sva_dfm_2, input_mem_banks_bank_a_50_sva_dfm_2,
          input_mem_banks_bank_a_51_sva_dfm_2, input_mem_banks_bank_a_52_sva_dfm_2,
          input_mem_banks_bank_a_53_sva_dfm_2, input_mem_banks_bank_a_54_sva_dfm_2,
          input_mem_banks_bank_a_55_sva_dfm_2, input_mem_banks_bank_a_56_sva_dfm_2,
          input_mem_banks_bank_a_57_sva_dfm_2, input_mem_banks_bank_a_58_sva_dfm_2,
          input_mem_banks_bank_a_59_sva_dfm_2, input_mem_banks_bank_a_60_sva_dfm_2,
          input_mem_banks_bank_a_61_sva_dfm_2, input_mem_banks_bank_a_62_sva_dfm_2,
          input_mem_banks_bank_a_63_sva_dfm_2, input_mem_banks_bank_a_64_sva_dfm_2,
          input_mem_banks_bank_a_65_sva_dfm_2, input_mem_banks_bank_a_66_sva_dfm_2,
          input_mem_banks_bank_a_67_sva_dfm_2, input_mem_banks_bank_a_68_sva_dfm_2,
          input_mem_banks_bank_a_69_sva_dfm_2, input_mem_banks_bank_a_70_sva_dfm_2,
          input_mem_banks_bank_a_71_sva_dfm_2, input_mem_banks_bank_a_72_sva_dfm_2,
          input_mem_banks_bank_a_73_sva_dfm_2, input_mem_banks_bank_a_74_sva_dfm_2,
          input_mem_banks_bank_a_75_sva_dfm_2, input_mem_banks_bank_a_76_sva_dfm_2,
          input_mem_banks_bank_a_77_sva_dfm_2, input_mem_banks_bank_a_78_sva_dfm_2,
          input_mem_banks_bank_a_79_sva_dfm_2, input_mem_banks_bank_a_80_sva_dfm_2,
          input_mem_banks_bank_a_81_sva_dfm_2, input_mem_banks_bank_a_82_sva_dfm_2,
          input_mem_banks_bank_a_83_sva_dfm_2, input_mem_banks_bank_a_84_sva_dfm_2,
          input_mem_banks_bank_a_85_sva_dfm_2, input_mem_banks_bank_a_86_sva_dfm_2,
          input_mem_banks_bank_a_87_sva_dfm_2, input_mem_banks_bank_a_88_sva_dfm_2,
          input_mem_banks_bank_a_89_sva_dfm_2, input_mem_banks_bank_a_90_sva_dfm_2,
          input_mem_banks_bank_a_91_sva_dfm_2, input_mem_banks_bank_a_92_sva_dfm_2,
          input_mem_banks_bank_a_93_sva_dfm_2, input_mem_banks_bank_a_94_sva_dfm_2,
          input_mem_banks_bank_a_95_sva_dfm_2, input_mem_banks_bank_a_96_sva_dfm_2,
          input_mem_banks_bank_a_97_sva_dfm_2, input_mem_banks_bank_a_98_sva_dfm_2,
          input_mem_banks_bank_a_99_sva_dfm_2, input_mem_banks_bank_a_100_sva_dfm_2,
          input_mem_banks_bank_a_101_sva_dfm_2, input_mem_banks_bank_a_102_sva_dfm_2,
          input_mem_banks_bank_a_103_sva_dfm_2, input_mem_banks_bank_a_104_sva_dfm_2,
          input_mem_banks_bank_a_105_sva_dfm_2, input_mem_banks_bank_a_106_sva_dfm_2,
          input_mem_banks_bank_a_107_sva_dfm_2, input_mem_banks_bank_a_108_sva_dfm_2,
          input_mem_banks_bank_a_109_sva_dfm_2, input_mem_banks_bank_a_110_sva_dfm_2,
          input_mem_banks_bank_a_111_sva_dfm_2, input_mem_banks_bank_a_112_sva_dfm_2,
          input_mem_banks_bank_a_113_sva_dfm_2, input_mem_banks_bank_a_114_sva_dfm_2,
          input_mem_banks_bank_a_115_sva_dfm_2, input_mem_banks_bank_a_116_sva_dfm_2,
          input_mem_banks_bank_a_117_sva_dfm_2, input_mem_banks_bank_a_118_sva_dfm_2,
          input_mem_banks_bank_a_119_sva_dfm_2, input_mem_banks_bank_a_120_sva_dfm_2,
          input_mem_banks_bank_a_121_sva_dfm_2, input_mem_banks_bank_a_122_sva_dfm_2,
          input_mem_banks_bank_a_123_sva_dfm_2, input_mem_banks_bank_a_124_sva_dfm_2,
          input_mem_banks_bank_a_125_sva_dfm_2, input_mem_banks_bank_a_126_sva_dfm_2,
          input_mem_banks_bank_a_127_sva_dfm_2, input_mem_banks_bank_a_128_sva_dfm_2,
          input_mem_banks_bank_a_129_sva_dfm_2, input_mem_banks_bank_a_130_sva_dfm_2,
          input_mem_banks_bank_a_131_sva_dfm_2, input_mem_banks_bank_a_132_sva_dfm_2,
          input_mem_banks_bank_a_133_sva_dfm_2, input_mem_banks_bank_a_134_sva_dfm_2,
          input_mem_banks_bank_a_135_sva_dfm_2, input_mem_banks_bank_a_136_sva_dfm_2,
          input_mem_banks_bank_a_137_sva_dfm_2, input_mem_banks_bank_a_138_sva_dfm_2,
          input_mem_banks_bank_a_139_sva_dfm_2, input_mem_banks_bank_a_140_sva_dfm_2,
          input_mem_banks_bank_a_141_sva_dfm_2, input_mem_banks_bank_a_142_sva_dfm_2,
          input_mem_banks_bank_a_143_sva_dfm_2, input_mem_banks_bank_a_144_sva_dfm_2,
          input_mem_banks_bank_a_145_sva_dfm_2, input_mem_banks_bank_a_146_sva_dfm_2,
          input_mem_banks_bank_a_147_sva_dfm_2, input_mem_banks_bank_a_148_sva_dfm_2,
          input_mem_banks_bank_a_149_sva_dfm_2, input_mem_banks_bank_a_150_sva_dfm_2,
          input_mem_banks_bank_a_151_sva_dfm_2, input_mem_banks_bank_a_152_sva_dfm_2,
          input_mem_banks_bank_a_153_sva_dfm_2, input_mem_banks_bank_a_154_sva_dfm_2,
          input_mem_banks_bank_a_155_sva_dfm_2, input_mem_banks_bank_a_156_sva_dfm_2,
          input_mem_banks_bank_a_157_sva_dfm_2, input_mem_banks_bank_a_158_sva_dfm_2,
          input_mem_banks_bank_a_159_sva_dfm_2, input_mem_banks_bank_a_160_sva_dfm_2,
          input_mem_banks_bank_a_161_sva_dfm_2, input_mem_banks_bank_a_162_sva_dfm_2,
          input_mem_banks_bank_a_163_sva_dfm_2, input_mem_banks_bank_a_164_sva_dfm_2,
          input_mem_banks_bank_a_165_sva_dfm_2, input_mem_banks_bank_a_166_sva_dfm_2,
          input_mem_banks_bank_a_167_sva_dfm_2, input_mem_banks_bank_a_168_sva_dfm_2,
          input_mem_banks_bank_a_169_sva_dfm_2, input_mem_banks_bank_a_170_sva_dfm_2,
          input_mem_banks_bank_a_171_sva_dfm_2, input_mem_banks_bank_a_172_sva_dfm_2,
          input_mem_banks_bank_a_173_sva_dfm_2, input_mem_banks_bank_a_174_sva_dfm_2,
          input_mem_banks_bank_a_175_sva_dfm_2, input_mem_banks_bank_a_176_sva_dfm_2,
          input_mem_banks_bank_a_177_sva_dfm_2, input_mem_banks_bank_a_178_sva_dfm_2,
          input_mem_banks_bank_a_179_sva_dfm_2, input_mem_banks_bank_a_180_sva_dfm_2,
          input_mem_banks_bank_a_181_sva_dfm_2, input_mem_banks_bank_a_182_sva_dfm_2,
          input_mem_banks_bank_a_183_sva_dfm_2, input_mem_banks_bank_a_184_sva_dfm_2,
          input_mem_banks_bank_a_185_sva_dfm_2, input_mem_banks_bank_a_186_sva_dfm_2,
          input_mem_banks_bank_a_187_sva_dfm_2, input_mem_banks_bank_a_188_sva_dfm_2,
          input_mem_banks_bank_a_189_sva_dfm_2, input_mem_banks_bank_a_190_sva_dfm_2,
          input_mem_banks_bank_a_191_sva_dfm_2, input_mem_banks_bank_a_192_sva_dfm_2,
          input_mem_banks_bank_a_193_sva_dfm_2, input_mem_banks_bank_a_194_sva_dfm_2,
          input_mem_banks_bank_a_195_sva_dfm_2, input_mem_banks_bank_a_196_sva_dfm_2,
          input_mem_banks_bank_a_197_sva_dfm_2, input_mem_banks_bank_a_198_sva_dfm_2,
          input_mem_banks_bank_a_199_sva_dfm_2, input_mem_banks_bank_a_200_sva_dfm_2,
          input_mem_banks_bank_a_201_sva_dfm_2, input_mem_banks_bank_a_202_sva_dfm_2,
          input_mem_banks_bank_a_203_sva_dfm_2, input_mem_banks_bank_a_204_sva_dfm_2,
          input_mem_banks_bank_a_205_sva_dfm_2, input_mem_banks_bank_a_206_sva_dfm_2,
          input_mem_banks_bank_a_207_sva_dfm_2, input_mem_banks_bank_a_208_sva_dfm_2,
          input_mem_banks_bank_a_209_sva_dfm_2, input_mem_banks_bank_a_210_sva_dfm_2,
          input_mem_banks_bank_a_211_sva_dfm_2, input_mem_banks_bank_a_212_sva_dfm_2,
          input_mem_banks_bank_a_213_sva_dfm_2, input_mem_banks_bank_a_214_sva_dfm_2,
          input_mem_banks_bank_a_215_sva_dfm_2, input_mem_banks_bank_a_216_sva_dfm_2,
          input_mem_banks_bank_a_217_sva_dfm_2, input_mem_banks_bank_a_218_sva_dfm_2,
          input_mem_banks_bank_a_219_sva_dfm_2, input_mem_banks_bank_a_220_sva_dfm_2,
          input_mem_banks_bank_a_221_sva_dfm_2, input_mem_banks_bank_a_222_sva_dfm_2,
          input_mem_banks_bank_a_223_sva_dfm_2, input_mem_banks_bank_a_224_sva_dfm_2,
          input_mem_banks_bank_a_225_sva_dfm_2, input_mem_banks_bank_a_226_sva_dfm_2,
          input_mem_banks_bank_a_227_sva_dfm_2, input_mem_banks_bank_a_228_sva_dfm_2,
          input_mem_banks_bank_a_229_sva_dfm_2, input_mem_banks_bank_a_230_sva_dfm_2,
          input_mem_banks_bank_a_231_sva_dfm_2, input_mem_banks_bank_a_232_sva_dfm_2,
          input_mem_banks_bank_a_233_sva_dfm_2, input_mem_banks_bank_a_234_sva_dfm_2,
          input_mem_banks_bank_a_235_sva_dfm_2, input_mem_banks_bank_a_236_sva_dfm_2,
          input_mem_banks_bank_a_237_sva_dfm_2, input_mem_banks_bank_a_238_sva_dfm_2,
          input_mem_banks_bank_a_239_sva_dfm_2, input_mem_banks_bank_a_240_sva_dfm_2,
          input_mem_banks_bank_a_241_sva_dfm_2, input_mem_banks_bank_a_242_sva_dfm_2,
          input_mem_banks_bank_a_243_sva_dfm_2, input_mem_banks_bank_a_244_sva_dfm_2,
          input_mem_banks_bank_a_245_sva_dfm_2, input_mem_banks_bank_a_246_sva_dfm_2,
          input_mem_banks_bank_a_247_sva_dfm_2, input_mem_banks_bank_a_248_sva_dfm_2,
          input_mem_banks_bank_a_249_sva_dfm_2, input_mem_banks_bank_a_250_sva_dfm_2,
          input_mem_banks_bank_a_251_sva_dfm_2, input_mem_banks_bank_a_252_sva_dfm_2,
          input_mem_banks_bank_a_253_sva_dfm_2, input_mem_banks_bank_a_254_sva_dfm_2,
          input_mem_banks_bank_a_255_sva_dfm_2, input_mem_banks_read_1_for_mux_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( input_read_req_valid_and_3_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= input_read_req_valid_lpi_1_dfm_1_6;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_15_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_146_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= rva_out_reg_data_30_25_sva_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_147_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= rva_out_reg_data_23_17_sva_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_7 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_148_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_7 <= rva_out_reg_data_15_9_sva_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_149_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= rva_out_reg_data_35_32_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_150_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_2 <= rva_out_reg_data_39_36_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_151_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2 <= rva_out_reg_data_46_40_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_4_2 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_152_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_4_2 <= rva_out_reg_data_62_48_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_153_enex5 ) begin
      rva_out_reg_data_127_112_sva_dfm_4_2 <= rva_out_reg_data_127_112_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_96_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_154_enex5 ) begin
      rva_out_reg_data_111_96_sva_dfm_4_2 <= rva_out_reg_data_111_96_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_80_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_155_enex5 ) begin
      rva_out_reg_data_95_80_sva_dfm_4_2 <= rva_out_reg_data_95_80_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_156_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_4_2 <= rva_out_reg_data_79_64_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_114_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_114_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_118_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_118_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_122_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_122_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_126_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_126_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_130_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_130_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_134_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_134_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_138_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_138_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_142_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_142_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_146_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_146_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_150_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_150_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_154_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_154_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_158_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_158_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_162_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_162_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_166_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_166_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_170_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_170_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_174_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_174_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_178_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_178_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_182_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_182_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_186_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_186_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_190_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_190_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_194_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_194_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_198_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_198_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_202_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_202_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_206_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_206_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_210_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_210_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_214_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_214_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_218_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_218_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_222_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_222_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_226_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_226_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_230_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_230_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_234_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_234_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_238_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_238_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_242_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_242_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_246_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_246_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_250_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_250_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_254_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_254_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_258_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_258_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_262_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_262_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_266_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_266_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_270_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_270_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_274_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_274_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_278_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_278_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_282_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_282_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_286_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_286_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_290_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_290_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_294_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_294_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_298_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_298_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_302_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_302_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_306_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_306_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_310_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_310_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_314_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_314_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_318_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_318_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_322_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_322_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_326_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_326_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_330_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_330_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_334_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_334_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_338_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_338_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_342_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_342_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_346_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_346_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_350_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_350_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_354_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_354_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_358_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_358_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_362_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_362_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_366_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_366_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_370_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_370_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_374_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_374_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_378_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_378_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_382_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_382_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_386_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_386_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_390_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_390_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_394_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_394_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_398_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_398_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_402_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_402_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_406_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_406_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_410_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_410_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_414_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_414_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_418_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_418_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_422_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_422_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_426_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_426_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_430_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_430_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_434_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_434_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_438_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_438_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_442_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_442_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_446_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_446_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_450_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_450_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_454_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_454_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_458_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_458_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_462_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_462_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_466_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_466_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_470_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_470_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_474_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_474_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_478_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_478_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_482_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_482_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_486_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_486_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_490_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_490_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_494_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_494_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_498_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_498_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_502_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_502_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_506_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_506_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_510_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_510_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_514_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_514_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_518_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_518_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_522_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_522_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_526_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_526_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_530_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_530_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_534_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_534_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_538_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_538_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_542_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_542_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_546_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_546_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_550_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_550_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_554_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_554_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_558_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_558_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_562_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_562_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_566_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_566_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_570_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_570_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_574_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_574_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_578_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_578_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_582_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_582_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_586_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_586_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_590_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_590_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_594_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_594_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_598_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_598_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_602_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_602_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_606_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_606_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_610_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_610_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_614_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_614_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_618_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_618_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_622_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_622_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_626_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_626_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_630_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_630_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_634_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_634_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_638_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_638_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_642_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_642_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_646_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_646_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_650_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_650_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_654_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_654_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_658_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_658_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_662_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_662_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_666_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_666_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_670_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_670_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_674_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_674_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_678_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_678_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_682_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_682_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_686_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_686_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_690_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_690_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_694_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_694_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_698_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_698_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_702_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_702_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_706_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_706_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_710_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_710_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_714_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_714_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_718_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_718_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_722_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_722_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_726_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_726_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_730_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_730_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_734_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_734_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_738_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_738_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_742_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_742_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_746_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_746_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_750_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_750_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_754_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_754_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_758_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_758_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_762_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_762_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_766_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_766_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_770_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_770_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_774_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_774_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_778_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_778_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_782_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_782_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_786_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_786_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_790_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_790_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_794_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_794_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_798_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_798_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_802_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_802_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_806_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_806_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_810_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_810_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_814_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_814_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_818_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_818_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_822_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_822_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_826_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_826_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_830_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_830_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_834_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_834_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_838_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_838_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_842_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_842_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_846_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_846_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_850_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_850_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_854_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_854_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_858_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_858_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_862_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_862_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_866_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_866_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_870_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_870_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_874_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_874_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_878_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_878_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_882_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_882_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_886_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_886_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_890_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_890_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_894_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_894_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_898_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_898_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_902_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_902_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_906_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_906_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_910_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_910_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_914_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_914_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_918_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_918_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_922_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_922_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_926_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_926_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_930_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_930_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_934_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_934_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_938_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_938_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_942_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_942_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_946_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_946_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_950_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_950_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_954_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_954_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_958_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_958_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_962_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_962_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_966_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_966_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_970_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_970_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_974_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_974_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_978_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_978_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_982_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_982_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_986_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_986_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_990_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_990_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_994_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_994_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_998_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_998_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1002_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1002_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1006_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1006_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1010_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1010_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1014_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1014_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1018_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1018_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1022_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1022_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1026_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1026_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1030_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1030_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1034_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1034_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1038_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1038_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1042_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1042_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1046_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1046_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1050_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1050_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1054_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1054_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1058_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1058_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1062_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1062_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1066_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1066_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1070_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1070_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1074_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1074_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1078_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1078_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1082_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1082_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1086_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1086_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1090_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1090_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1094_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1094_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1098_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1098_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1102_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1102_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1106_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1106_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1110_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1110_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1114_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1114_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1118_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1118_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1122_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1122_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1126_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1126_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1130_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1130_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1134_rgt) & while_stage_0_3 ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= MUX_v_128_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1134_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_86_nl) & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_6 <= 1'b0;
      rva_in_reg_rw_sva_st_6 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_15_cse ) begin
      rva_in_reg_rw_sva_st_1_6 <= rva_in_reg_rw_sva_st_1_5;
      rva_in_reg_rw_sva_st_6 <= rva_in_reg_rw_sva_st_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_36_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_4[0];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_4[8];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[16];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[31];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_64_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_65_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:9];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_66_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:17];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_67_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[30:25];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( input_read_req_valid_and_4_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_9_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_19_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_4 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_157_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_4 <= rva_out_reg_data_30_25_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_158_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_4 <= rva_out_reg_data_23_17_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_6 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_159_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_6 <= rva_out_reg_data_15_9_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= 4'b0000;
      rva_out_reg_data_39_36_sva_dfm_4_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_4_1 <= 7'b0000000;
      rva_out_reg_data_62_48_sva_dfm_4_1 <= 15'b000000000000000;
    end
    else if ( and_1235_cse ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= MUX1HOT_v_4_4_2(rva_out_reg_data_35_32_sva_dfm_1_5,
          rva_out_reg_data_35_32_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[35:32]),
          (weight_port_read_out_data_0_2_sva_dfm_mx0w1_14_0[3:0]), {PECore_PushAxiRsp_if_asn_69
          , PECore_PushAxiRsp_if_asn_71 , PECore_PushAxiRsp_if_asn_67 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_39_36_sva_dfm_4_1 <= MUX1HOT_v_4_4_2(rva_out_reg_data_39_36_sva_dfm_1_5,
          rva_out_reg_data_39_36_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:36]),
          (weight_port_read_out_data_0_2_sva_dfm_mx0w1_14_0[7:4]), {PECore_PushAxiRsp_if_asn_69
          , PECore_PushAxiRsp_if_asn_71 , PECore_PushAxiRsp_if_asn_67 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_46_40_sva_dfm_4_1 <= MUX1HOT_v_7_4_2(rva_out_reg_data_46_40_sva_dfm_1_5,
          rva_out_reg_data_46_40_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[46:40]),
          (weight_port_read_out_data_0_2_sva_dfm_mx0w1_14_0[14:8]), {PECore_PushAxiRsp_if_asn_69
          , PECore_PushAxiRsp_if_asn_71 , PECore_PushAxiRsp_if_asn_67 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_62_48_sva_dfm_4_1 <= MUX1HOT_v_15_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_14_0,
          rva_out_reg_data_62_48_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[62:48]),
          weight_port_read_out_data_0_3_sva_dfm_mx0w3_14_0, {PECore_PushAxiRsp_if_asn_69
          , PECore_PushAxiRsp_if_asn_71 , PECore_PushAxiRsp_if_asn_67 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_111_96_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_95_80_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_79_64_sva_dfm_4_1 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_72_cse ) begin
      rva_out_reg_data_127_112_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_127_112_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000003,
          weight_port_read_out_data_1_3_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_665 , and_dcpl_666});
      rva_out_reg_data_111_96_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_111_96_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000002,
          weight_port_read_out_data_1_2_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_665 , and_dcpl_666});
      rva_out_reg_data_95_80_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_95_80_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000005,
          weight_port_read_out_data_1_5_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_665 , and_dcpl_666});
      rva_out_reg_data_79_64_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_79_64_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_15_0_000004,
          weight_port_read_out_data_1_4_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_665 , and_dcpl_666});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_6 <= 15'b000000000000000;
      rva_out_reg_data_46_40_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_39_36_sva_dfm_6 <= 4'b0000;
      rva_out_reg_data_35_32_sva_dfm_6 <= 4'b0000;
    end
    else if ( and_1252_cse ) begin
      rva_out_reg_data_62_48_sva_dfm_6 <= rva_out_reg_data_62_48_sva_dfm_6_mx1;
      rva_out_reg_data_46_40_sva_dfm_6 <= rva_out_reg_data_46_40_sva_dfm_6_mx1;
      rva_out_reg_data_39_36_sva_dfm_6 <= rva_out_reg_data_39_36_sva_dfm_6_mx1;
      rva_out_reg_data_35_32_sva_dfm_6 <= rva_out_reg_data_35_32_sva_dfm_6_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_18_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & ((and_dcpl_212 & rva_in_reg_rw_sva_5) | PECore_PushAxiRsp_mux_18_itm_1_mx0c1)
        ) begin
      PECore_PushAxiRsp_mux_18_itm_1 <= MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
          weight_port_read_out_data_mux_18_nl, PECore_PushAxiRsp_mux_18_itm_1_mx0c1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~(while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5))
        | rva_in_reg_rw_sva_5)) ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          weight_port_read_out_data_0_2_sva_dfm_mx0w1_15, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_45_tmp ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= MUX1HOT_v_128_3_2(input_mem_banks_read_read_data_lpi_1_dfm_1_3,
          weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d, weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1,
          {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          , and_676_nl , nor_383_nl});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_160_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_5 <= rva_out_reg_data_46_40_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_5 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_161_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_5 <= rva_out_reg_data_39_36_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_5 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_162_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_5 <= rva_out_reg_data_35_32_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_95_80_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_111_96_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_127_112_sva_dfm_6 <= 16'b0000000000000000;
    end
    else if ( and_1272_cse ) begin
      rva_out_reg_data_79_64_sva_dfm_6 <= rva_out_reg_data_79_64_sva_dfm_4_mx0w0;
      rva_out_reg_data_95_80_sva_dfm_6 <= rva_out_reg_data_95_80_sva_dfm_4_mx0w0;
      rva_out_reg_data_111_96_sva_dfm_6 <= rva_out_reg_data_111_96_sva_dfm_4_mx0w0;
      rva_out_reg_data_127_112_sva_dfm_6 <= rva_out_reg_data_127_112_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_5
          <= 1'b0;
    end
    else if ( rva_out_reg_data_and_80_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_base_input_and_tmp ) begin
      pe_manager_base_input_sva <= MUX_v_15_2_2(pe_manager_base_input_sva_dfm_3_1,
          PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl,
          and_dcpl_197);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( (~((~((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6:4]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:7]!=3'b000))) & nor_438_cse
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:12]!=3'b000))) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]))
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) & rva_in_PopNB_mioi_return_rsc_z_mxwt
        & nor_472_cse & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18:17]==2'b10) &
        rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)) & while_stage_0_3)) & rva_in_reg_rw_and_4_cse
        ) begin
      pe_manager_base_input_sva_dfm_3_1 <= MUX_v_15_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[62:48]),
          pe_manager_base_input_sva_mx1, or_422_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_21_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_23_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= MUX_s_1_2_2(weight_mem_run_3_for_5_and_158_nl,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= MUX_s_1_2_2(weight_mem_run_3_for_5_and_151_nl,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= MUX_s_1_2_2(weight_mem_run_3_for_5_and_100_nl,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= MUX_s_1_2_2(weight_mem_run_3_for_5_and_112_nl,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_3 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_163_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_3 <= rva_out_reg_data_30_25_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_164_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_3 <= rva_out_reg_data_23_17_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_165_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_5 <= rva_out_reg_data_15_9_sva_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_26_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_3 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_46_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_27_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_nl,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_166_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= rva_out_reg_data_30_25_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_167_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= rva_out_reg_data_23_17_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_168_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= rva_out_reg_data_15_9_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_169_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= rva_out_reg_data_35_32_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_170_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= rva_out_reg_data_39_36_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_171_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= rva_out_reg_data_46_40_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_1_4 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_172_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_1_4 <= rva_out_reg_data_62_48_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]))) & while_stage_0_4 )
        begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_31_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_47_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ reg_rva_in_reg_rw_sva_2_cse) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= input_read_req_valid_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= 6'b000000;
      rva_out_reg_data_23_17_sva_dfm_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_97_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= MUX_v_6_2_2(6'b000000, (pe_manager_base_weight_sva_mx2[14:9]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
      rva_out_reg_data_23_17_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_base_weight_sva_mx2[7:1]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_173_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= rva_out_reg_data_15_9_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_174_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= rva_out_reg_data_35_32_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_175_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= rva_out_reg_data_39_36_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_176_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= rva_out_reg_data_46_40_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_1_3 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_177_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_1_3 <= rva_out_reg_data_62_48_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_35_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_36_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_104_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= rva_out_reg_data_15_9_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_178_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= rva_out_reg_data_35_32_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_179_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= rva_out_reg_data_39_36_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_180_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= rva_out_reg_data_46_40_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_1_2 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_181_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_1_2 <= pe_manager_base_input_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (and_dcpl_481 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        & while_stage_0_3 ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_2_1,
          PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_481 & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1==4'b0100)
        & and_dcpl_488 & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3))
        & and_dcpl_189 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_40_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ reg_rva_in_reg_rw_sva_st_1_1_cse) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
        & while_stage_0_3 ) begin
      input_read_req_valid_lpi_1_dfm_1_2 <= input_read_req_valid_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_1 <= 7'b0000000;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3;
      rva_out_reg_data_15_9_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_num_input_sva[7:1]),
          and_289_cse);
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_45_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_1 <= pe_config_is_cluster_sva;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= pe_config_is_bias_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (or_dcpl_132 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
        | (~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))))
        & and_dcpl_197 ) begin
      input_read_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= 1'b0;
      rva_out_reg_data_35_32_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_39_36_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_1_1 <= 7'b0000000;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_49_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= (pe_config_num_output_sva[7]) & (~(and_289_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1))
          & PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
      rva_out_reg_data_35_32_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl
          & (signext_4_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1)) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_39_36_sva_dfm_1_1 <= (pe_manager_base_bias_sva[7:4]) & ({{3{and_289_cse}},
          and_289_cse}) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_46_40_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl
          & (signext_7_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1)) & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_15 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(mux_2_itm & (~((~ rva_in_reg_rw_sva_st_1_5) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3))
        & while_stage_0_6)) & and_dcpl_212 ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_15 <= mux1h_1_nl & (~ or_dcpl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_14_0 <= 15'b000000000000000;
    end
    else if ( and_1313_tmp ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_14_0 <= MUX_v_15_2_2(15'b000000000000000,
          mux1h_7_nl, not_1918_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_15
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_14_0
          <= 15'b000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_25_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_15
          <= weight_mem_banks_load_store_for_else_mux1h_28_nl & (~ or_dcpl_309);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_14_0
          <= MUX_v_15_2_2(15'b000000000000000, weight_mem_banks_load_store_for_else_mux1h_44_nl,
          not_1861_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_2_15_1 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_76_cse ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_0 <= weight_port_read_out_data_0_1_sva_dfm_1_15;
      weight_port_read_out_data_0_0_sva_dfm_2_15_1 <= weight_port_read_out_data_0_0_sva_dfm_1_1_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_88_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_1 <= weight_port_read_out_data_0_1_sva_dfm_1_14_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_5_rsp_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_89_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_5_rsp_1 <= weight_port_read_out_data_0_1_sva_dfm_4_14_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_1_14_0 <= 15'b000000000000000;
    end
    else if ( mux_342_nl & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & while_stage_0_7 & PECoreRun_wen ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_1_14_0 <= MUX1HOT_v_15_9_2(weight_port_read_out_data_0_1_sva_mx0_14_0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[30:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[30:16]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[30:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[30:16]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[30:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[30:16]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[30:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[14:0]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55
          , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_179_cse , weight_mem_run_3_for_5_and_180_ssc
          , weight_mem_run_3_for_5_and_181_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_4_14_0 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_90_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_4_14_0 <= reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_15
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_72_nl) ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_15
          <= mux1h_3_nl & (~ mux_259_tmp);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_14_0
          <= 15'b000000000000000;
    end
    else if ( (~ mux_350_nl) & PECoreRun_wen ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_14_0
          <= MUX_v_15_2_2(15'b000000000000000, mux1h_8_nl, not_1920_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_1_15 <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_1_1_14_0 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_63_ssc ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_1_15 <= MUX_s_1_2_2(weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_15,
          weight_port_read_out_data_0_0_sva_dfm_mx0w1_15, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
      weight_port_read_out_data_0_0_sva_dfm_1_1_14_0 <= MUX_v_15_2_2(weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_14_0,
          weight_port_read_out_data_0_0_sva_dfm_mx0w1_14_0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1_14_0 <= 15'b000000000000000;
    end
    else if ( mux_354_nl & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & while_stage_0_7 & PECoreRun_wen ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1_14_0 <= MUX1HOT_v_15_9_2(weight_port_read_out_data_0_3_sva_mx0_14_0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[62:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[62:48]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[62:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[62:48]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[62:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[62:48]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[62:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[46:32]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_55
          , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse
          , weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse
          , weight_mem_run_3_for_5_and_195_ssc , weight_mem_run_3_for_5_and_188_cse
          , weight_mem_run_3_for_5_and_181_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_15 <= 1'b0;
    end
    else if ( PECoreRun_wen & (and_dcpl_212 | and_dcpl_48) ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_15 <= MUX_s_1_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w1_15,
          weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_15, and_dcpl_48);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_14_0 <= 15'b000000000000000;
    end
    else if ( mux_357_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_14_0 <= MUX_v_15_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w1_14_0,
          weight_port_read_out_data_0_0_sva_dfm_1_mx0w0_14_0, and_dcpl_48);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_15
          <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_84_nl ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_15
          <= MUX_s_1_2_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl,
          weight_port_read_out_data_0_2_sva_dfm_mx0w1_15, or_dcpl_277);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0
          <= 15'b000000000000000;
    end
    else if ( mux_363_nl & PECoreRun_wen ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0
          <= MUX_v_15_2_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_64_nl,
          weight_port_read_out_data_0_2_sva_dfm_mx0w1_14_0, or_dcpl_277);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_91_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1 <= weight_port_read_out_data_0_0_sva_dfm_2_14_0_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_14_0_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_92_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_14_0_1 <= weight_port_read_out_data_0_0_sva_dfm_1_1_14_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_126_enex5 | rva_out_reg_data_and_113_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_enexo <= rva_out_reg_data_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_125_enex5 | rva_out_reg_data_and_114_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_enexo <= rva_out_reg_data_and_125_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_124_enex5 | rva_out_reg_data_and_115_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_7_enexo <= rva_out_reg_data_and_124_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_131_enex5 | rva_out_reg_data_and_116_enex5 ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_4_enexo <= rva_out_reg_data_and_131_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_132_enex5 | rva_out_reg_data_and_117_enex5 ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_4_enexo <= rva_out_reg_data_and_132_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_133_enex5 | rva_out_reg_data_and_118_enex5 ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_4_enexo <= rva_out_reg_data_and_133_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_enex5 | rva_out_reg_data_and_119_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_4_enexo <= rva_out_reg_data_and_134_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_130_enex5 | rva_out_reg_data_and_120_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_4_enexo <= rva_out_reg_data_and_130_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_129_enex5 | rva_out_reg_data_and_121_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo <= rva_out_reg_data_and_129_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_128_enex5 | rva_out_reg_data_and_122_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_enexo <= rva_out_reg_data_and_128_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_127_enex5 | rva_out_reg_data_and_123_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo <= rva_out_reg_data_and_127_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_86_enex5 | weight_port_read_out_data_and_78_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_4_1_enexo <= weight_port_read_out_data_and_86_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_52_enex5 | input_mem_banks_read_read_data_and_48_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo
          <= input_mem_banks_read_read_data_and_52_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_53_enex5 | input_mem_banks_read_read_data_and_49_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo
          <= input_mem_banks_read_read_data_and_53_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_54_enex5 | input_mem_banks_read_read_data_and_50_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo
          <= input_mem_banks_read_read_data_and_54_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_55_enex5 | input_mem_banks_read_read_data_and_51_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo
          <= input_mem_banks_read_read_data_and_55_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_1_enex5 | input_mem_banks_read_1_read_data_and_5_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_1_read_data_and_1_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp | weight_port_read_out_data_and_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000000
          <= data_in_tmp_operator_2_for_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_79_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000000
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000001
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_80_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000001
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000002
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_81_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000002
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000003
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_82_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000003
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000004
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_83_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000004
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000005
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_84_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000005
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000006
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_85_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_128_127_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_16_1000006
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_2_enex5 | input_mem_banks_read_1_read_data_and_1_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= input_mem_banks_read_1_read_data_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( weight_read_addrs_and_5_cse | weight_read_addrs_and_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= weight_read_addrs_and_5_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_6_14_1_lpi_1_dfm_1_enexo <= 1'b1;
    end
    else if ( weight_read_addrs_and_7_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_weight_read_addrs_6_14_1_lpi_1_dfm_1_enexo <= weight_read_addrs_and_7_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= 1'b1;
    end
    else if ( weight_read_addrs_and_5_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= weight_read_addrs_and_5_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_6_14_1_lpi_1_dfm_1_enexo_1 <= 1'b1;
    end
    else if ( weight_read_addrs_and_7_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_read_addrs_6_14_1_lpi_1_dfm_1_enexo_1 <= weight_read_addrs_and_7_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= 1'b1;
    end
    else if ( operator_15_false_1_and_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= operator_15_false_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= 1'b1;
    end
    else if ( weight_read_addrs_and_5_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= weight_read_addrs_and_5_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo_1
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo_1
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_32_enex5 | weight_write_data_data_and_24_enex5
        ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_32_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_33_enex5 | weight_write_data_data_and_25_enex5
        ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_33_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_34_enex5 | weight_write_data_data_and_26_enex5
        ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_34_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_35_enex5 | weight_write_data_data_and_27_enex5
        ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_35_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_36_enex5 | weight_write_data_data_and_28_enex5
        ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_36_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_37_enex5 | weight_write_data_data_and_29_enex5
        ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_37_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_38_enex5 | weight_write_data_data_and_30_enex5
        ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_38_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_39_enex5 | weight_write_data_data_and_31_enex5
        ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_39_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_write_addrs_and_3_enex5 | weight_write_addrs_and_enex5 ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= weight_write_addrs_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_32_enex5 ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_33_enex5 ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_34_enex5 ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_35_enex5 ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_36_enex5 ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_37_enex5 ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_38_enex5 ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_39_enex5 ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_addrs_and_3_enex5 ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_read_addrs_and_29_enex5 ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_config_num_output_enexo <= 1'b1;
    end
    else if ( pe_config_num_manager_and_cse | pe_config_UpdateManagerCounter_if_if_and_enex5
        ) begin
      reg_pe_config_num_output_enexo <= pe_config_num_manager_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_read_addrs_and_30_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_data_sva_1_enexo <= 1'b1;
    end
    else if ( rva_in_reg_data_and_tmp | PEManager_15U_PEManagerWrite_and_enex5 )
        begin
      reg_rva_in_reg_data_sva_1_enexo <= rva_in_reg_data_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_56_enex5 | input_mem_banks_read_read_data_and_52_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo
          <= input_mem_banks_read_read_data_and_56_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_57_enex5 | input_mem_banks_read_read_data_and_53_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo
          <= input_mem_banks_read_read_data_and_57_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_58_enex5 | input_mem_banks_read_read_data_and_54_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo
          <= input_mem_banks_read_read_data_and_58_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_59_enex5 | input_mem_banks_read_read_data_and_55_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo
          <= input_mem_banks_read_read_data_and_59_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 | input_mem_banks_read_1_read_data_and_2_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_1_read_data_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_135_enex5 | rva_out_reg_data_and_124_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= rva_out_reg_data_and_135_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_136_enex5 | rva_out_reg_data_and_125_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= rva_out_reg_data_and_136_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_137_enex5 | rva_out_reg_data_and_126_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= rva_out_reg_data_and_137_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_91_enex5 | weight_port_read_out_data_and_86_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_91_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_138_enex5 | rva_out_reg_data_and_127_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= rva_out_reg_data_and_138_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_139_enex5 | rva_out_reg_data_and_128_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo <= rva_out_reg_data_and_139_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_140_enex5 | rva_out_reg_data_and_129_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo <= rva_out_reg_data_and_140_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_141_enex5 | rva_out_reg_data_and_130_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_3_enexo <= rva_out_reg_data_and_141_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_142_enex5 | rva_out_reg_data_and_131_enex5 ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_3_enexo <= rva_out_reg_data_and_142_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_143_enex5 | rva_out_reg_data_and_132_enex5 ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_3_enexo <= rva_out_reg_data_and_143_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_144_enex5 | rva_out_reg_data_and_133_enex5 ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_3_enexo <= rva_out_reg_data_and_144_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_145_enex5 | rva_out_reg_data_and_134_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_3_enexo <= rva_out_reg_data_and_145_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_60_enex5 | input_mem_banks_read_read_data_and_56_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= input_mem_banks_read_read_data_and_60_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_61_enex5 | input_mem_banks_read_read_data_and_57_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= input_mem_banks_read_read_data_and_61_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_62_enex5 | input_mem_banks_read_read_data_and_58_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= input_mem_banks_read_read_data_and_62_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_63_enex5 | input_mem_banks_read_read_data_and_59_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= input_mem_banks_read_read_data_and_63_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp | input_mem_banks_read_1_read_data_and_3_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= input_mem_banks_read_1_read_data_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_146_enex5 | rva_out_reg_data_and_135_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= rva_out_reg_data_and_146_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_147_enex5 | rva_out_reg_data_and_136_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= rva_out_reg_data_and_147_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_148_enex5 | rva_out_reg_data_and_137_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= rva_out_reg_data_and_148_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_88_enex5 | weight_port_read_out_data_and_87_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_88_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_149_enex5 | rva_out_reg_data_and_138_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= rva_out_reg_data_and_149_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_150_enex5 | rva_out_reg_data_and_139_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo <= rva_out_reg_data_and_150_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_151_enex5 | rva_out_reg_data_and_140_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo <= rva_out_reg_data_and_151_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_152_enex5 | rva_out_reg_data_and_141_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_2_enexo <= rva_out_reg_data_and_152_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_153_enex5 | rva_out_reg_data_and_142_enex5 ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_2_enexo <= rva_out_reg_data_and_153_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_154_enex5 | rva_out_reg_data_and_143_enex5 ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_2_enexo <= rva_out_reg_data_and_154_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_155_enex5 | rva_out_reg_data_and_144_enex5 ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_2_enexo <= rva_out_reg_data_and_155_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_156_enex5 | rva_out_reg_data_and_145_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_2_enexo <= rva_out_reg_data_and_156_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= 1'b1;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_1_for_and_cse | weight_mem_write_arbxbar_xbar_for_empty_and_enex5
        ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= weight_mem_write_arbxbar_xbar_for_1_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_64_enex5 | input_mem_banks_read_read_data_and_60_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= input_mem_banks_read_read_data_and_64_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_65_enex5 | input_mem_banks_read_read_data_and_61_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo
          <= input_mem_banks_read_read_data_and_65_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_66_enex5 | input_mem_banks_read_read_data_and_62_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= input_mem_banks_read_read_data_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_67_enex5 | input_mem_banks_read_read_data_and_63_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= input_mem_banks_read_read_data_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_157_enex5 | rva_out_reg_data_and_146_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_4_enexo <= rva_out_reg_data_and_157_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_158_enex5 | rva_out_reg_data_and_147_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_4_enexo <= rva_out_reg_data_and_158_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_159_enex5 | rva_out_reg_data_and_148_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_6_enexo <= rva_out_reg_data_and_159_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1235_cse | rva_out_reg_data_and_149_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= and_1235_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1235_cse | rva_out_reg_data_and_150_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo <= and_1235_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1235_cse | rva_out_reg_data_and_151_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo <= and_1235_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1235_cse | rva_out_reg_data_and_152_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_1_enexo <= and_1235_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_72_cse | rva_out_reg_data_and_153_enex5 ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_1_enexo <= rva_out_reg_data_and_72_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_72_cse | rva_out_reg_data_and_154_enex5 ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_1_enexo <= rva_out_reg_data_and_72_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_72_cse | rva_out_reg_data_and_155_enex5 ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_1_enexo <= rva_out_reg_data_and_72_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_72_cse | rva_out_reg_data_and_156_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_1_enexo <= rva_out_reg_data_and_72_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_45_tmp | input_mem_banks_read_read_data_and_64_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_read_data_and_45_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_45_tmp | input_mem_banks_read_read_data_and_65_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1 <= input_mem_banks_read_read_data_and_45_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_45_tmp | input_mem_banks_read_read_data_and_66_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2 <= input_mem_banks_read_read_data_and_45_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_3 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_45_tmp | input_mem_banks_read_read_data_and_67_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_3 <= input_mem_banks_read_read_data_and_45_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_163_enex5 | rva_out_reg_data_and_157_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_3_enexo <= rva_out_reg_data_and_163_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_164_enex5 | rva_out_reg_data_and_158_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_3_enexo <= rva_out_reg_data_and_164_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_165_enex5 | rva_out_reg_data_and_159_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_5_enexo <= rva_out_reg_data_and_165_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_171_enex5 | rva_out_reg_data_and_160_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_4_enexo <= rva_out_reg_data_and_171_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_170_enex5 | rva_out_reg_data_and_161_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_4_enexo <= rva_out_reg_data_and_170_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_169_enex5 | rva_out_reg_data_and_162_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_4_enexo <= rva_out_reg_data_and_169_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_166_enex5 | rva_out_reg_data_and_163_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_2_enexo <= rva_out_reg_data_and_166_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_167_enex5 | rva_out_reg_data_and_164_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_2_enexo <= rva_out_reg_data_and_167_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_168_enex5 | rva_out_reg_data_and_165_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_4_enexo <= rva_out_reg_data_and_168_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_47_enex5 | input_mem_banks_read_read_data_and_46_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_read_data_and_47_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_97_cse | rva_out_reg_data_and_166_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= rva_out_reg_data_and_97_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_97_cse | rva_out_reg_data_and_167_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= rva_out_reg_data_and_97_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_173_enex5 | rva_out_reg_data_and_168_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= rva_out_reg_data_and_173_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_174_enex5 | rva_out_reg_data_and_169_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= rva_out_reg_data_and_174_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_175_enex5 | rva_out_reg_data_and_170_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= rva_out_reg_data_and_175_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_176_enex5 | rva_out_reg_data_and_171_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= rva_out_reg_data_and_176_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_177_enex5 | rva_out_reg_data_and_172_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_1_3_enexo <= rva_out_reg_data_and_177_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp | input_mem_banks_read_read_data_and_47_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1 <= input_mem_banks_read_1_read_data_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_104_enex5 | rva_out_reg_data_and_173_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= rva_out_reg_data_and_104_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_178_enex5 | rva_out_reg_data_and_174_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= rva_out_reg_data_and_178_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_179_enex5 | rva_out_reg_data_and_175_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= rva_out_reg_data_and_179_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_180_enex5 | rva_out_reg_data_and_176_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= rva_out_reg_data_and_180_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_181_enex5 | rva_out_reg_data_and_177_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_1_2_enexo <= rva_out_reg_data_and_181_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse | rva_out_reg_data_and_104_enex5
        ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_49_cse | rva_out_reg_data_and_178_enex5
        ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_49_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_49_cse | rva_out_reg_data_and_179_enex5
        ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_49_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_49_cse | rva_out_reg_data_and_180_enex5
        ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_49_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_input_enexo <= 1'b1;
    end
    else if ( pe_manager_base_input_and_tmp | rva_out_reg_data_and_181_enex5 ) begin
      reg_pe_manager_base_input_enexo <= pe_manager_base_input_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1313_tmp | weight_port_read_out_data_and_88_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo <= and_1313_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_90_enex5 | weight_port_read_out_data_and_89_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_4_1_enexo <= weight_port_read_out_data_and_90_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_87_enex5 | weight_port_read_out_data_and_90_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_87_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_92_enex5 | weight_port_read_out_data_and_91_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_92_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_63_ssc | weight_port_read_out_data_and_92_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_1_enexo <= weight_port_read_out_data_and_63_ssc;
    end
  end
  assign nl_operator_4_false_acc_nl = pe_config_manager_counter_sva_mx1 + 4'b0001;
  assign operator_4_false_acc_nl = nl_operator_4_false_acc_nl[3:0];
  assign pe_config_UpdateManagerCounter_if_not_7_nl = ~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  assign nl_input_read_addrs_sva_1_1  = pe_config_input_counter_sva_mx1 + (pe_manager_base_input_sva_mx1[7:0]);
  assign PECore_UpdateFSM_switch_lp_not_27_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_not_28_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_not_29_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_not_30_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_not_31_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_not_19_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign nl_ProductSum_for_acc_14_itm_1  = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_5_cmp_31_z);
  assign mux_286_nl = MUX_s_1_2_2(not_tmp_469, mux_tmp_268, or_691_cse);
  assign mux_285_nl = MUX_s_1_2_2(not_tmp_469, mux_tmp_268, or_687_cse);
  assign mux_287_nl = MUX_s_1_2_2(mux_286_nl, mux_285_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_127_16_mx0[111:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign or_771_nl = (weight_read_addrs_5_lpi_1_dfm_3_2_0[1:0]!=2'b00);
  assign mux_306_nl = MUX_s_1_2_2((~ (weight_read_addrs_5_lpi_1_dfm_3_2_0[1])), (weight_read_addrs_5_lpi_1_dfm_3_2_0[1]),
      weight_read_addrs_5_lpi_1_dfm_3_2_0[0]);
  assign mux_307_nl = MUX_s_1_2_2(or_771_nl, mux_306_nl, weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign mux_308_nl = MUX_s_1_2_2((weight_read_addrs_3_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_3_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_3_lpi_1_dfm_3_2_0[0]);
  assign mux_309_nl = MUX_s_1_2_2(mux_308_nl, nor_428_cse, weight_read_addrs_3_lpi_1_dfm_3_2_0[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_76_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[15:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_76_nl);
  assign nor_264_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_4_nl = MUX_s_1_2_2(nor_264_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_72_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[15:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_72_nl);
  assign nor_265_nl = ~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_5_nl = MUX_s_1_2_2(nor_265_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_54_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_22_nl = (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp);
  assign or_20_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_6_nl = MUX_s_1_2_2(or_22_nl, or_20_nl, while_stage_0_6);
  assign or_27_nl = (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6])))
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign or_25_nl = (~(Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6 |
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3))
      | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_7_nl = MUX_s_1_2_2(or_25_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3,
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1);
  assign mux_8_nl = MUX_s_1_2_2(or_27_nl, mux_7_nl, while_stage_0_5);
  assign or_23_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_9_nl = MUX_s_1_2_2(mux_8_nl, or_23_nl, while_stage_0_6);
  assign mux_10_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_3, (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign nor_429_nl = ~((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign nor_430_nl = ~((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | (~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | (~ reg_rva_in_reg_rw_sva_st_1_1_cse));
  assign mux_310_nl = MUX_s_1_2_2(nor_429_nl, nor_430_nl, while_stage_0_3);
  assign mux_311_nl = MUX_s_1_2_2(mux_310_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2,
      while_stage_0_4);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl
      = MUX_v_11_2_2(11'b00000000000, PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign mux_312_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_5_1, nor_431_cse,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl = (state_mux_1_cse!=2'b00)
      | state_0_sva_mx1;
  assign PECore_UpdateFSM_switch_lp_or_nl = PECore_UpdateFSM_switch_lp_equal_tmp_6
      | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  assign PECore_UpdateFSM_switch_lp_mux1h_15_nl = MUX1HOT_v_2_3_2((signext_2_1(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl)),
      2'b01, 2'b10, {PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      , PECore_UpdateFSM_switch_lp_or_nl , PECore_RunScale_PECore_RunScale_if_and_1_svs_1});
  assign PECore_UpdateFSM_switch_lp_nor_8_nl = ~(PECore_PushOutput_PECore_PushOutput_if_and_svs_1
      | PECore_UpdateFSM_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_and_1_nl = MUX_v_2_2_2(2'b00, PECore_UpdateFSM_switch_lp_mux1h_15_nl,
      PECore_UpdateFSM_switch_lp_nor_8_nl);
  assign mux_313_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_3_1, nor_431_cse,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_314_nl = MUX_s_1_2_2(and_1331_cse, nor_431_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nl_operator_8_false_acc_sdt_sva_1  = conv_u2s_8_9(pe_config_num_output_sva)
      + 9'b111111111;
  assign PECore_UpdateFSM_switch_lp_not_38_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_not_21_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign mux_35_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_4_lpi_1_dfm_1, (~ rva_in_reg_rw_sva_st_1_4),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_2_nl
      = ~((weight_read_addrs_1_lpi_1_dfm_2_2_0!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl = (weight_read_addrs_1_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_20_nl = (weight_read_addrs_1_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_nl = (weight_read_addrs_1_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_24_nl = (weight_read_addrs_1_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign or_180_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ or_dcpl_59);
  assign mux_36_nl = MUX_s_1_2_2(or_dcpl_63, or_180_nl, while_stage_0_5);
  assign or_181_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ or_dcpl_52);
  assign mux_37_nl = MUX_s_1_2_2(or_dcpl_64, or_181_nl, while_stage_0_5);
  assign or_184_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 | and_739_cse));
  assign mux_38_nl = MUX_s_1_2_2(or_187_cse, or_184_nl, while_stage_0_5);
  assign mux_373_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp,
      and_733_cse, weight_mem_read_arbxbar_xbar_1_for_3_1_operator_7_false_1_operator_7_false_1_or_tmp);
  assign mux_46_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp,
      mux_373_nl, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign mux_45_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp,
      and_733_cse, and_740_cse);
  assign mux_47_nl = MUX_s_1_2_2(mux_46_nl, mux_45_nl, Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7);
  assign mux_48_nl = MUX_s_1_2_2(mux_47_nl, mux_tmp_44, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]);
  assign mux_49_nl = MUX_s_1_2_2(mux_48_nl, mux_256_cse, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign mux_50_nl = MUX_s_1_2_2(mux_49_nl, mux_tmp_44, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign mux_51_nl = MUX_s_1_2_2(mux_50_nl, mux_256_cse, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign mux_52_nl = MUX_s_1_2_2(mux_51_nl, mux_tmp_42, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign mux_53_nl = MUX_s_1_2_2(mux_52_nl, mux_256_cse, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign mux_39_nl = MUX_s_1_2_2(and_741_cse, and_742_cse, nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_tmp);
  assign mux_43_nl = MUX_s_1_2_2(mux_tmp_42, mux_39_nl, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1);
  assign mux_54_nl = MUX_s_1_2_2(mux_53_nl, mux_43_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign or_201_nl = (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ mux_54_nl);
  assign or_190_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ or_dcpl_31);
  assign mux_55_nl = MUX_s_1_2_2(or_201_nl, or_190_nl, while_stage_0_5);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl
      = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]), pe_config_is_zero_first_sva_mx1,
      PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_19_nl
      = MUX_s_1_2_2(PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl,
      pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_or_5_cse_1);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_129_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_101_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_115_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_122_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_94_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_108_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_130_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_102_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_116_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_123_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_95_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_109_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_131_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_103_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_117_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_124_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_96_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_110_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_132_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_104_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_118_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_125_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_97_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_111_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_133_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign and_938_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])
      & (~ or_639_tmp);
  assign and_939_nl = and_dcpl_643 & (~ or_639_tmp);
  assign and_940_nl = nor_275_cse & (~ or_639_tmp);
  assign mux1h_2_nl = MUX1HOT_v_16_3_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[63:48]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[63:48]), (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[31:16]),
      {and_938_nl , and_939_nl , and_940_nl});
  assign not_1864_nl = ~ or_639_tmp;
  assign mux_62_nl = MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]),
      (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_63_nl = MUX_s_1_2_2(mux_62_nl, nor_275_cse, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_126_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_127_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_128_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_112_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_114_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign and_658_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign and_660_nl = and_dcpl_652 & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign and_664_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      & and_dcpl_655;
  assign and_668_nl = (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      & weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_669_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_load_store_for_else_mux1h_37_nl = MUX1HOT_v_16_5_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[47:32]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[47:32]), (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[15:0]),
      (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[15:0]), (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[15:0]),
      {and_658_nl , and_660_nl , and_664_nl , and_668_nl , and_669_nl});
  assign and_661_nl = and_dcpl_652 & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]));
  assign weight_mem_banks_load_store_for_else_or_nl = MUX_v_16_2_2(weight_mem_banks_load_store_for_else_mux1h_37_nl,
      16'b1111111111111111, and_661_nl);
  assign or_643_nl = ((~((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]) | (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2])))
      & and_dcpl_652) | (and_dcpl_655 & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_275_nl = MUX_v_16_2_2(weight_mem_banks_load_store_for_else_or_nl, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[15:0]),
      or_643_nl);
  assign nor_398_nl = ~((mux_tmp_256 & and_dcpl_652) | (and_dcpl_724 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4));
  assign mux_79_nl = MUX_s_1_2_2(or_tmp_67, (~ mux_tmp_76), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_78_nl = MUX_s_1_2_2((~ mux_tmp_76), or_tmp_67, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_80_nl = MUX_s_1_2_2(mux_79_nl, mux_78_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_77_nl = MUX_s_1_2_2((~ mux_tmp_76), or_tmp_67, or_202_cse);
  assign mux_81_nl = MUX_s_1_2_2(mux_80_nl, mux_77_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_113_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_78_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b110)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b011)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_38_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b101)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_nl = (pe_manager_base_weight_sva[1])
      & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_133_itm_1 & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_nl = (pe_manager_base_weight_sva[2])
      & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_145_itm_1 & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_5_itm_1
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_nl = (pe_manager_base_weight_sva[2])
      & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_4_itm_1
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign mux_85_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, (~ pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_973_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & fsm_output;
  assign input_mem_banks_read_1_for_mux_nl = MUX_v_8_2_2(input_read_addrs_sva_1_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4,
      and_973_nl);
  assign mux_86_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign weight_port_read_out_data_mux_18_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_18_mx0w2,
      weight_port_read_out_data_0_3_sva_dfm_mx0w3_15, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_676_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign nor_383_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl
      = pe_manager_base_input_sva_mx1 & ({{14{and_289_cse}}, and_289_cse}) & ({{14{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
  assign or_422_nl = or_dcpl_132 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) |
      (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | or_dcpl_273;
  assign weight_mem_run_3_for_5_and_158_nl = (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_lpi_1_dfm_1;
  assign weight_mem_run_3_for_5_and_151_nl = (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_lpi_1_dfm_1;
  assign weight_mem_run_3_for_5_and_100_nl = (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_lpi_1_dfm_1;
  assign weight_mem_run_3_for_5_and_112_nl = (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_nl = (pe_manager_base_weight_sva[1:0]==2'b11)
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1 & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_2,
      (pe_manager_base_weight_sva_mx1_3_0[0]), PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2,
      (pe_manager_base_weight_sva_mx2[8]), PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl =
      (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl = MUX_s_1_2_2(pe_config_is_valid_sva,
      pe_manager_zero_active_sva, and_289_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl = MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1,
      (pe_manager_num_input_sva[0]), and_289_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl = MUX_v_4_2_2(pe_config_num_manager_sva,
      (pe_manager_base_bias_sva[3:0]), and_289_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl = MUX_v_7_2_2((pe_config_num_output_sva[6:0]),
      (pe_manager_base_bias_sva[14:8]), and_289_cse);
  assign mux1h_1_nl = MUX1HOT_s_1_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_15,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1[15]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_15,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1[15]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1[15]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[31]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[31]),
      weight_port_read_out_data_0_1_sva_mx0_15, {and_929_cse , and_930_cse , and_931_cse
      , and_932_cse , and_933_cse , and_934_cse , and_935_cse , nor_397_cse});
  assign mux1h_7_nl = MUX1HOT_v_15_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1[14:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_14_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1[14:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1[14:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[30:16]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[30:16]),
      weight_port_read_out_data_0_1_sva_mx0_14_0, {and_929_cse , and_930_cse , and_931_cse
      , and_932_cse , and_933_cse , and_934_cse , and_935_cse , nor_397_cse});
  assign not_1918_nl = ~ or_dcpl;
  assign weight_mem_banks_load_store_for_else_mux1h_28_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[63]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[31]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[31]),
      {and_647_ssc , and_648_ssc , and_649_ssc});
  assign weight_mem_banks_load_store_for_else_mux1h_44_nl = MUX1HOT_v_15_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[62:48]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[30:16]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[30:16]),
      rva_out_reg_data_62_48_sva_dfm_1_4, {and_647_ssc , and_648_ssc , and_649_ssc
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_1861_nl = ~ or_dcpl_309;
  assign mux_341_nl = MUX_s_1_2_2(not_tmp_653, mux_tmp_323, or_691_cse);
  assign mux_340_nl = MUX_s_1_2_2(not_tmp_653, mux_tmp_323, or_687_cse);
  assign mux_342_nl = MUX_s_1_2_2(mux_341_nl, mux_340_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux1h_3_nl = MUX1HOT_s_1_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[47]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[15]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[15]),
      weight_port_read_out_data_0_3_sva_dfm_mx0w3_15, {and_654_ssc , and_656_ssc
      , and_657_ssc , or_dcpl_277});
  assign mux_70_nl = MUX_s_1_2_2(mux_tmp_65, (~ mux_tmp_67), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_69_nl = MUX_s_1_2_2((~ mux_tmp_67), mux_tmp_65, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_71_nl = MUX_s_1_2_2(mux_70_nl, mux_69_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_68_nl = MUX_s_1_2_2((~ mux_tmp_67), mux_tmp_65, or_202_cse);
  assign mux_72_nl = MUX_s_1_2_2(mux_71_nl, mux_68_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign mux1h_8_nl = MUX1HOT_v_15_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[46:32]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[14:0]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[14:0]),
      weight_port_read_out_data_0_3_sva_dfm_mx0w3_14_0, {and_654_ssc , and_656_ssc
      , and_657_ssc , or_dcpl_277});
  assign not_1920_nl = ~ mux_259_tmp;
  assign or_903_nl = weight_mem_run_3_for_land_1_lpi_1_dfm_2 | not_tmp_658;
  assign mux_343_nl = MUX_s_1_2_2((~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])),
      (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_344_nl = MUX_s_1_2_2(mux_343_nl, or_202_cse, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign mux_348_nl = MUX_s_1_2_2(not_tmp_658, mux_344_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_349_nl = MUX_s_1_2_2(or_903_nl, mux_348_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_350_nl = MUX_s_1_2_2(not_tmp_658, mux_349_nl, while_stage_0_6);
  assign mux_353_nl = MUX_s_1_2_2(not_tmp_662, mux_tmp_335, or_691_cse);
  assign mux_352_nl = MUX_s_1_2_2(not_tmp_662, mux_tmp_335, or_687_cse);
  assign mux_354_nl = MUX_s_1_2_2(mux_353_nl, mux_352_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_916_nl = reg_weight_mem_run_3_for_5_and_168_itm_2_cse | reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_166_itm_2_cse | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | weight_mem_run_3_for_5_and_164_itm_2 | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_162_itm_2_cse | and_1339_cse;
  assign and_1340_nl = ((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[1])
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_2)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign and_1341_nl = ((~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[1]))
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_2)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign mux_355_nl = MUX_s_1_2_2(and_1340_nl, and_1341_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[2]);
  assign and_1342_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_2)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign mux_356_nl = MUX_s_1_2_2(mux_355_nl, and_1342_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_3[0]);
  assign or_914_nl = or_tmp_425 | mux_356_nl;
  assign mux_357_nl = MUX_s_1_2_2(or_916_nl, or_914_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl
      = (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[31]) & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]));
  assign mux_82_nl = MUX_s_1_2_2((~ or_tmp_59), or_tmp_61, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1);
  assign mux_83_nl = MUX_s_1_2_2((~ or_tmp_60), mux_82_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_84_nl = MUX_s_1_2_2(and_dcpl_212, mux_83_nl, while_stage_0_6);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_136_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_64_nl
      = MUX_v_15_2_2(15'b000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[30:16]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_136_nl);
  assign nor_477_nl = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_2 | (~ and_tmp_24));
  assign mux_361_nl = MUX_s_1_2_2(and_tmp_24, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_362_nl = MUX_s_1_2_2(nor_477_nl, mux_361_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_363_nl = MUX_s_1_2_2(and_tmp_24, mux_362_nl, while_stage_0_6);

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_6_2;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [5:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_9_2;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [8:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_8_2;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [7:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    result = result | (input_5 & {11{sel[5]}});
    result = result | (input_6 & {11{sel[6]}});
    result = result | (input_7 & {11{sel[7]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function automatic [127:0] MUX1HOT_v_128_3_2;
    input [127:0] input_2;
    input [127:0] input_1;
    input [127:0] input_0;
    input [2:0] sel;
    reg [127:0] result;
  begin
    result = input_0 & {128{sel[0]}};
    result = result | (input_1 & {128{sel[1]}});
    result = result | (input_2 & {128{sel[2]}});
    MUX1HOT_v_128_3_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_3_2;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [2:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | (input_1 & {15{sel[1]}});
    result = result | (input_2 & {15{sel[2]}});
    MUX1HOT_v_15_3_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_4_2;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [3:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | (input_1 & {15{sel[1]}});
    result = result | (input_2 & {15{sel[2]}});
    result = result | (input_3 & {15{sel[3]}});
    MUX1HOT_v_15_4_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_8_2;
    input [14:0] input_7;
    input [14:0] input_6;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [7:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | (input_1 & {15{sel[1]}});
    result = result | (input_2 & {15{sel[2]}});
    result = result | (input_3 & {15{sel[3]}});
    result = result | (input_4 & {15{sel[4]}});
    result = result | (input_5 & {15{sel[5]}});
    result = result | (input_6 & {15{sel[6]}});
    result = result | (input_7 & {15{sel[7]}});
    MUX1HOT_v_15_8_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_9_2;
    input [14:0] input_8;
    input [14:0] input_7;
    input [14:0] input_6;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [8:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | (input_1 & {15{sel[1]}});
    result = result | (input_2 & {15{sel[2]}});
    result = result | (input_3 & {15{sel[3]}});
    result = result | (input_4 & {15{sel[4]}});
    result = result | (input_5 & {15{sel[5]}});
    result = result | (input_6 & {15{sel[6]}});
    result = result | (input_7 & {15{sel[7]}});
    result = result | (input_8 & {15{sel[8]}});
    MUX1HOT_v_15_9_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_5_2;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [4:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    MUX1HOT_v_16_5_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_6_2;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [5:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    MUX1HOT_v_16_6_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_8_2;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [7:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    result = result | (input_7 & {16{sel[7]}});
    MUX1HOT_v_16_8_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_9_2;
    input [15:0] input_8;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [8:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    result = result | (input_7 & {16{sel[7]}});
    result = result | (input_8 & {16{sel[8]}});
    MUX1HOT_v_16_9_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | (input_1 & {32{sel[1]}});
    result = result | (input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_8_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input [2:0] sel;
    reg  result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_s_1_8_2 = result;
  end
  endfunction


  function automatic [111:0] MUX_v_112_2_2;
    input [111:0] input_0;
    input [111:0] input_1;
    input  sel;
    reg [111:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_112_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_8_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [10:0] input_2;
    input [10:0] input_3;
    input [10:0] input_4;
    input [10:0] input_5;
    input [10:0] input_6;
    input [10:0] input_7;
    input [2:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_11_8_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_256_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [127:0] input_2;
    input [127:0] input_3;
    input [127:0] input_4;
    input [127:0] input_5;
    input [127:0] input_6;
    input [127:0] input_7;
    input [127:0] input_8;
    input [127:0] input_9;
    input [127:0] input_10;
    input [127:0] input_11;
    input [127:0] input_12;
    input [127:0] input_13;
    input [127:0] input_14;
    input [127:0] input_15;
    input [127:0] input_16;
    input [127:0] input_17;
    input [127:0] input_18;
    input [127:0] input_19;
    input [127:0] input_20;
    input [127:0] input_21;
    input [127:0] input_22;
    input [127:0] input_23;
    input [127:0] input_24;
    input [127:0] input_25;
    input [127:0] input_26;
    input [127:0] input_27;
    input [127:0] input_28;
    input [127:0] input_29;
    input [127:0] input_30;
    input [127:0] input_31;
    input [127:0] input_32;
    input [127:0] input_33;
    input [127:0] input_34;
    input [127:0] input_35;
    input [127:0] input_36;
    input [127:0] input_37;
    input [127:0] input_38;
    input [127:0] input_39;
    input [127:0] input_40;
    input [127:0] input_41;
    input [127:0] input_42;
    input [127:0] input_43;
    input [127:0] input_44;
    input [127:0] input_45;
    input [127:0] input_46;
    input [127:0] input_47;
    input [127:0] input_48;
    input [127:0] input_49;
    input [127:0] input_50;
    input [127:0] input_51;
    input [127:0] input_52;
    input [127:0] input_53;
    input [127:0] input_54;
    input [127:0] input_55;
    input [127:0] input_56;
    input [127:0] input_57;
    input [127:0] input_58;
    input [127:0] input_59;
    input [127:0] input_60;
    input [127:0] input_61;
    input [127:0] input_62;
    input [127:0] input_63;
    input [127:0] input_64;
    input [127:0] input_65;
    input [127:0] input_66;
    input [127:0] input_67;
    input [127:0] input_68;
    input [127:0] input_69;
    input [127:0] input_70;
    input [127:0] input_71;
    input [127:0] input_72;
    input [127:0] input_73;
    input [127:0] input_74;
    input [127:0] input_75;
    input [127:0] input_76;
    input [127:0] input_77;
    input [127:0] input_78;
    input [127:0] input_79;
    input [127:0] input_80;
    input [127:0] input_81;
    input [127:0] input_82;
    input [127:0] input_83;
    input [127:0] input_84;
    input [127:0] input_85;
    input [127:0] input_86;
    input [127:0] input_87;
    input [127:0] input_88;
    input [127:0] input_89;
    input [127:0] input_90;
    input [127:0] input_91;
    input [127:0] input_92;
    input [127:0] input_93;
    input [127:0] input_94;
    input [127:0] input_95;
    input [127:0] input_96;
    input [127:0] input_97;
    input [127:0] input_98;
    input [127:0] input_99;
    input [127:0] input_100;
    input [127:0] input_101;
    input [127:0] input_102;
    input [127:0] input_103;
    input [127:0] input_104;
    input [127:0] input_105;
    input [127:0] input_106;
    input [127:0] input_107;
    input [127:0] input_108;
    input [127:0] input_109;
    input [127:0] input_110;
    input [127:0] input_111;
    input [127:0] input_112;
    input [127:0] input_113;
    input [127:0] input_114;
    input [127:0] input_115;
    input [127:0] input_116;
    input [127:0] input_117;
    input [127:0] input_118;
    input [127:0] input_119;
    input [127:0] input_120;
    input [127:0] input_121;
    input [127:0] input_122;
    input [127:0] input_123;
    input [127:0] input_124;
    input [127:0] input_125;
    input [127:0] input_126;
    input [127:0] input_127;
    input [127:0] input_128;
    input [127:0] input_129;
    input [127:0] input_130;
    input [127:0] input_131;
    input [127:0] input_132;
    input [127:0] input_133;
    input [127:0] input_134;
    input [127:0] input_135;
    input [127:0] input_136;
    input [127:0] input_137;
    input [127:0] input_138;
    input [127:0] input_139;
    input [127:0] input_140;
    input [127:0] input_141;
    input [127:0] input_142;
    input [127:0] input_143;
    input [127:0] input_144;
    input [127:0] input_145;
    input [127:0] input_146;
    input [127:0] input_147;
    input [127:0] input_148;
    input [127:0] input_149;
    input [127:0] input_150;
    input [127:0] input_151;
    input [127:0] input_152;
    input [127:0] input_153;
    input [127:0] input_154;
    input [127:0] input_155;
    input [127:0] input_156;
    input [127:0] input_157;
    input [127:0] input_158;
    input [127:0] input_159;
    input [127:0] input_160;
    input [127:0] input_161;
    input [127:0] input_162;
    input [127:0] input_163;
    input [127:0] input_164;
    input [127:0] input_165;
    input [127:0] input_166;
    input [127:0] input_167;
    input [127:0] input_168;
    input [127:0] input_169;
    input [127:0] input_170;
    input [127:0] input_171;
    input [127:0] input_172;
    input [127:0] input_173;
    input [127:0] input_174;
    input [127:0] input_175;
    input [127:0] input_176;
    input [127:0] input_177;
    input [127:0] input_178;
    input [127:0] input_179;
    input [127:0] input_180;
    input [127:0] input_181;
    input [127:0] input_182;
    input [127:0] input_183;
    input [127:0] input_184;
    input [127:0] input_185;
    input [127:0] input_186;
    input [127:0] input_187;
    input [127:0] input_188;
    input [127:0] input_189;
    input [127:0] input_190;
    input [127:0] input_191;
    input [127:0] input_192;
    input [127:0] input_193;
    input [127:0] input_194;
    input [127:0] input_195;
    input [127:0] input_196;
    input [127:0] input_197;
    input [127:0] input_198;
    input [127:0] input_199;
    input [127:0] input_200;
    input [127:0] input_201;
    input [127:0] input_202;
    input [127:0] input_203;
    input [127:0] input_204;
    input [127:0] input_205;
    input [127:0] input_206;
    input [127:0] input_207;
    input [127:0] input_208;
    input [127:0] input_209;
    input [127:0] input_210;
    input [127:0] input_211;
    input [127:0] input_212;
    input [127:0] input_213;
    input [127:0] input_214;
    input [127:0] input_215;
    input [127:0] input_216;
    input [127:0] input_217;
    input [127:0] input_218;
    input [127:0] input_219;
    input [127:0] input_220;
    input [127:0] input_221;
    input [127:0] input_222;
    input [127:0] input_223;
    input [127:0] input_224;
    input [127:0] input_225;
    input [127:0] input_226;
    input [127:0] input_227;
    input [127:0] input_228;
    input [127:0] input_229;
    input [127:0] input_230;
    input [127:0] input_231;
    input [127:0] input_232;
    input [127:0] input_233;
    input [127:0] input_234;
    input [127:0] input_235;
    input [127:0] input_236;
    input [127:0] input_237;
    input [127:0] input_238;
    input [127:0] input_239;
    input [127:0] input_240;
    input [127:0] input_241;
    input [127:0] input_242;
    input [127:0] input_243;
    input [127:0] input_244;
    input [127:0] input_245;
    input [127:0] input_246;
    input [127:0] input_247;
    input [127:0] input_248;
    input [127:0] input_249;
    input [127:0] input_250;
    input [127:0] input_251;
    input [127:0] input_252;
    input [127:0] input_253;
    input [127:0] input_254;
    input [127:0] input_255;
    input [7:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      8'b00000000 : begin
        result = input_0;
      end
      8'b00000001 : begin
        result = input_1;
      end
      8'b00000010 : begin
        result = input_2;
      end
      8'b00000011 : begin
        result = input_3;
      end
      8'b00000100 : begin
        result = input_4;
      end
      8'b00000101 : begin
        result = input_5;
      end
      8'b00000110 : begin
        result = input_6;
      end
      8'b00000111 : begin
        result = input_7;
      end
      8'b00001000 : begin
        result = input_8;
      end
      8'b00001001 : begin
        result = input_9;
      end
      8'b00001010 : begin
        result = input_10;
      end
      8'b00001011 : begin
        result = input_11;
      end
      8'b00001100 : begin
        result = input_12;
      end
      8'b00001101 : begin
        result = input_13;
      end
      8'b00001110 : begin
        result = input_14;
      end
      8'b00001111 : begin
        result = input_15;
      end
      8'b00010000 : begin
        result = input_16;
      end
      8'b00010001 : begin
        result = input_17;
      end
      8'b00010010 : begin
        result = input_18;
      end
      8'b00010011 : begin
        result = input_19;
      end
      8'b00010100 : begin
        result = input_20;
      end
      8'b00010101 : begin
        result = input_21;
      end
      8'b00010110 : begin
        result = input_22;
      end
      8'b00010111 : begin
        result = input_23;
      end
      8'b00011000 : begin
        result = input_24;
      end
      8'b00011001 : begin
        result = input_25;
      end
      8'b00011010 : begin
        result = input_26;
      end
      8'b00011011 : begin
        result = input_27;
      end
      8'b00011100 : begin
        result = input_28;
      end
      8'b00011101 : begin
        result = input_29;
      end
      8'b00011110 : begin
        result = input_30;
      end
      8'b00011111 : begin
        result = input_31;
      end
      8'b00100000 : begin
        result = input_32;
      end
      8'b00100001 : begin
        result = input_33;
      end
      8'b00100010 : begin
        result = input_34;
      end
      8'b00100011 : begin
        result = input_35;
      end
      8'b00100100 : begin
        result = input_36;
      end
      8'b00100101 : begin
        result = input_37;
      end
      8'b00100110 : begin
        result = input_38;
      end
      8'b00100111 : begin
        result = input_39;
      end
      8'b00101000 : begin
        result = input_40;
      end
      8'b00101001 : begin
        result = input_41;
      end
      8'b00101010 : begin
        result = input_42;
      end
      8'b00101011 : begin
        result = input_43;
      end
      8'b00101100 : begin
        result = input_44;
      end
      8'b00101101 : begin
        result = input_45;
      end
      8'b00101110 : begin
        result = input_46;
      end
      8'b00101111 : begin
        result = input_47;
      end
      8'b00110000 : begin
        result = input_48;
      end
      8'b00110001 : begin
        result = input_49;
      end
      8'b00110010 : begin
        result = input_50;
      end
      8'b00110011 : begin
        result = input_51;
      end
      8'b00110100 : begin
        result = input_52;
      end
      8'b00110101 : begin
        result = input_53;
      end
      8'b00110110 : begin
        result = input_54;
      end
      8'b00110111 : begin
        result = input_55;
      end
      8'b00111000 : begin
        result = input_56;
      end
      8'b00111001 : begin
        result = input_57;
      end
      8'b00111010 : begin
        result = input_58;
      end
      8'b00111011 : begin
        result = input_59;
      end
      8'b00111100 : begin
        result = input_60;
      end
      8'b00111101 : begin
        result = input_61;
      end
      8'b00111110 : begin
        result = input_62;
      end
      8'b00111111 : begin
        result = input_63;
      end
      8'b01000000 : begin
        result = input_64;
      end
      8'b01000001 : begin
        result = input_65;
      end
      8'b01000010 : begin
        result = input_66;
      end
      8'b01000011 : begin
        result = input_67;
      end
      8'b01000100 : begin
        result = input_68;
      end
      8'b01000101 : begin
        result = input_69;
      end
      8'b01000110 : begin
        result = input_70;
      end
      8'b01000111 : begin
        result = input_71;
      end
      8'b01001000 : begin
        result = input_72;
      end
      8'b01001001 : begin
        result = input_73;
      end
      8'b01001010 : begin
        result = input_74;
      end
      8'b01001011 : begin
        result = input_75;
      end
      8'b01001100 : begin
        result = input_76;
      end
      8'b01001101 : begin
        result = input_77;
      end
      8'b01001110 : begin
        result = input_78;
      end
      8'b01001111 : begin
        result = input_79;
      end
      8'b01010000 : begin
        result = input_80;
      end
      8'b01010001 : begin
        result = input_81;
      end
      8'b01010010 : begin
        result = input_82;
      end
      8'b01010011 : begin
        result = input_83;
      end
      8'b01010100 : begin
        result = input_84;
      end
      8'b01010101 : begin
        result = input_85;
      end
      8'b01010110 : begin
        result = input_86;
      end
      8'b01010111 : begin
        result = input_87;
      end
      8'b01011000 : begin
        result = input_88;
      end
      8'b01011001 : begin
        result = input_89;
      end
      8'b01011010 : begin
        result = input_90;
      end
      8'b01011011 : begin
        result = input_91;
      end
      8'b01011100 : begin
        result = input_92;
      end
      8'b01011101 : begin
        result = input_93;
      end
      8'b01011110 : begin
        result = input_94;
      end
      8'b01011111 : begin
        result = input_95;
      end
      8'b01100000 : begin
        result = input_96;
      end
      8'b01100001 : begin
        result = input_97;
      end
      8'b01100010 : begin
        result = input_98;
      end
      8'b01100011 : begin
        result = input_99;
      end
      8'b01100100 : begin
        result = input_100;
      end
      8'b01100101 : begin
        result = input_101;
      end
      8'b01100110 : begin
        result = input_102;
      end
      8'b01100111 : begin
        result = input_103;
      end
      8'b01101000 : begin
        result = input_104;
      end
      8'b01101001 : begin
        result = input_105;
      end
      8'b01101010 : begin
        result = input_106;
      end
      8'b01101011 : begin
        result = input_107;
      end
      8'b01101100 : begin
        result = input_108;
      end
      8'b01101101 : begin
        result = input_109;
      end
      8'b01101110 : begin
        result = input_110;
      end
      8'b01101111 : begin
        result = input_111;
      end
      8'b01110000 : begin
        result = input_112;
      end
      8'b01110001 : begin
        result = input_113;
      end
      8'b01110010 : begin
        result = input_114;
      end
      8'b01110011 : begin
        result = input_115;
      end
      8'b01110100 : begin
        result = input_116;
      end
      8'b01110101 : begin
        result = input_117;
      end
      8'b01110110 : begin
        result = input_118;
      end
      8'b01110111 : begin
        result = input_119;
      end
      8'b01111000 : begin
        result = input_120;
      end
      8'b01111001 : begin
        result = input_121;
      end
      8'b01111010 : begin
        result = input_122;
      end
      8'b01111011 : begin
        result = input_123;
      end
      8'b01111100 : begin
        result = input_124;
      end
      8'b01111101 : begin
        result = input_125;
      end
      8'b01111110 : begin
        result = input_126;
      end
      8'b01111111 : begin
        result = input_127;
      end
      8'b10000000 : begin
        result = input_128;
      end
      8'b10000001 : begin
        result = input_129;
      end
      8'b10000010 : begin
        result = input_130;
      end
      8'b10000011 : begin
        result = input_131;
      end
      8'b10000100 : begin
        result = input_132;
      end
      8'b10000101 : begin
        result = input_133;
      end
      8'b10000110 : begin
        result = input_134;
      end
      8'b10000111 : begin
        result = input_135;
      end
      8'b10001000 : begin
        result = input_136;
      end
      8'b10001001 : begin
        result = input_137;
      end
      8'b10001010 : begin
        result = input_138;
      end
      8'b10001011 : begin
        result = input_139;
      end
      8'b10001100 : begin
        result = input_140;
      end
      8'b10001101 : begin
        result = input_141;
      end
      8'b10001110 : begin
        result = input_142;
      end
      8'b10001111 : begin
        result = input_143;
      end
      8'b10010000 : begin
        result = input_144;
      end
      8'b10010001 : begin
        result = input_145;
      end
      8'b10010010 : begin
        result = input_146;
      end
      8'b10010011 : begin
        result = input_147;
      end
      8'b10010100 : begin
        result = input_148;
      end
      8'b10010101 : begin
        result = input_149;
      end
      8'b10010110 : begin
        result = input_150;
      end
      8'b10010111 : begin
        result = input_151;
      end
      8'b10011000 : begin
        result = input_152;
      end
      8'b10011001 : begin
        result = input_153;
      end
      8'b10011010 : begin
        result = input_154;
      end
      8'b10011011 : begin
        result = input_155;
      end
      8'b10011100 : begin
        result = input_156;
      end
      8'b10011101 : begin
        result = input_157;
      end
      8'b10011110 : begin
        result = input_158;
      end
      8'b10011111 : begin
        result = input_159;
      end
      8'b10100000 : begin
        result = input_160;
      end
      8'b10100001 : begin
        result = input_161;
      end
      8'b10100010 : begin
        result = input_162;
      end
      8'b10100011 : begin
        result = input_163;
      end
      8'b10100100 : begin
        result = input_164;
      end
      8'b10100101 : begin
        result = input_165;
      end
      8'b10100110 : begin
        result = input_166;
      end
      8'b10100111 : begin
        result = input_167;
      end
      8'b10101000 : begin
        result = input_168;
      end
      8'b10101001 : begin
        result = input_169;
      end
      8'b10101010 : begin
        result = input_170;
      end
      8'b10101011 : begin
        result = input_171;
      end
      8'b10101100 : begin
        result = input_172;
      end
      8'b10101101 : begin
        result = input_173;
      end
      8'b10101110 : begin
        result = input_174;
      end
      8'b10101111 : begin
        result = input_175;
      end
      8'b10110000 : begin
        result = input_176;
      end
      8'b10110001 : begin
        result = input_177;
      end
      8'b10110010 : begin
        result = input_178;
      end
      8'b10110011 : begin
        result = input_179;
      end
      8'b10110100 : begin
        result = input_180;
      end
      8'b10110101 : begin
        result = input_181;
      end
      8'b10110110 : begin
        result = input_182;
      end
      8'b10110111 : begin
        result = input_183;
      end
      8'b10111000 : begin
        result = input_184;
      end
      8'b10111001 : begin
        result = input_185;
      end
      8'b10111010 : begin
        result = input_186;
      end
      8'b10111011 : begin
        result = input_187;
      end
      8'b10111100 : begin
        result = input_188;
      end
      8'b10111101 : begin
        result = input_189;
      end
      8'b10111110 : begin
        result = input_190;
      end
      8'b10111111 : begin
        result = input_191;
      end
      8'b11000000 : begin
        result = input_192;
      end
      8'b11000001 : begin
        result = input_193;
      end
      8'b11000010 : begin
        result = input_194;
      end
      8'b11000011 : begin
        result = input_195;
      end
      8'b11000100 : begin
        result = input_196;
      end
      8'b11000101 : begin
        result = input_197;
      end
      8'b11000110 : begin
        result = input_198;
      end
      8'b11000111 : begin
        result = input_199;
      end
      8'b11001000 : begin
        result = input_200;
      end
      8'b11001001 : begin
        result = input_201;
      end
      8'b11001010 : begin
        result = input_202;
      end
      8'b11001011 : begin
        result = input_203;
      end
      8'b11001100 : begin
        result = input_204;
      end
      8'b11001101 : begin
        result = input_205;
      end
      8'b11001110 : begin
        result = input_206;
      end
      8'b11001111 : begin
        result = input_207;
      end
      8'b11010000 : begin
        result = input_208;
      end
      8'b11010001 : begin
        result = input_209;
      end
      8'b11010010 : begin
        result = input_210;
      end
      8'b11010011 : begin
        result = input_211;
      end
      8'b11010100 : begin
        result = input_212;
      end
      8'b11010101 : begin
        result = input_213;
      end
      8'b11010110 : begin
        result = input_214;
      end
      8'b11010111 : begin
        result = input_215;
      end
      8'b11011000 : begin
        result = input_216;
      end
      8'b11011001 : begin
        result = input_217;
      end
      8'b11011010 : begin
        result = input_218;
      end
      8'b11011011 : begin
        result = input_219;
      end
      8'b11011100 : begin
        result = input_220;
      end
      8'b11011101 : begin
        result = input_221;
      end
      8'b11011110 : begin
        result = input_222;
      end
      8'b11011111 : begin
        result = input_223;
      end
      8'b11100000 : begin
        result = input_224;
      end
      8'b11100001 : begin
        result = input_225;
      end
      8'b11100010 : begin
        result = input_226;
      end
      8'b11100011 : begin
        result = input_227;
      end
      8'b11100100 : begin
        result = input_228;
      end
      8'b11100101 : begin
        result = input_229;
      end
      8'b11100110 : begin
        result = input_230;
      end
      8'b11100111 : begin
        result = input_231;
      end
      8'b11101000 : begin
        result = input_232;
      end
      8'b11101001 : begin
        result = input_233;
      end
      8'b11101010 : begin
        result = input_234;
      end
      8'b11101011 : begin
        result = input_235;
      end
      8'b11101100 : begin
        result = input_236;
      end
      8'b11101101 : begin
        result = input_237;
      end
      8'b11101110 : begin
        result = input_238;
      end
      8'b11101111 : begin
        result = input_239;
      end
      8'b11110000 : begin
        result = input_240;
      end
      8'b11110001 : begin
        result = input_241;
      end
      8'b11110010 : begin
        result = input_242;
      end
      8'b11110011 : begin
        result = input_243;
      end
      8'b11110100 : begin
        result = input_244;
      end
      8'b11110101 : begin
        result = input_245;
      end
      8'b11110110 : begin
        result = input_246;
      end
      8'b11110111 : begin
        result = input_247;
      end
      8'b11111000 : begin
        result = input_248;
      end
      8'b11111001 : begin
        result = input_249;
      end
      8'b11111010 : begin
        result = input_250;
      end
      8'b11111011 : begin
        result = input_251;
      end
      8'b11111100 : begin
        result = input_252;
      end
      8'b11111101 : begin
        result = input_253;
      end
      8'b11111110 : begin
        result = input_254;
      end
      default : begin
        result = input_255;
      end
    endcase
    MUX_v_128_256_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input  sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input  sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_8_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [2:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_16_8_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [34:0] MUX_v_35_2_2;
    input [34:0] input_0;
    input [34:0] input_1;
    input  sel;
    reg [34:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_35_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [10:0] signext_11_1;
    input  vector;
  begin
    signext_11_1= {{10{vector}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input  vector;
  begin
    signext_4_1= {{3{vector}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input  vector;
  begin
    signext_7_1= {{6{vector}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [34:0] conv_u2u_34_35 ;
    input [33:0]  vector ;
  begin
    conv_u2u_34_35 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore
// ------------------------------------------------------------------


module PECore (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [137:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [168:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [127:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_c;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_en;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_c;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_5_en;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_z;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_clken;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_we;
  wire [127:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_1 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_1_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_1_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_1_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_2 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_2_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_2_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_2_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_3 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_3_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_3_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_3_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_4 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_4_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_4_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_4_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_5 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_5_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_5_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_5_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_6 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_6_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_6_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_6_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_7 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_7_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_7_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_7_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_8 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_8_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_8_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_8_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_9 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_9_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_9_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_9_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_10 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_10_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_10_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_10_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_11 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_11_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_11_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_11_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_12 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_12_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_12_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_12_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_13 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_13_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_13_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_13_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_14 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_14_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_14_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_14_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_15 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_15_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_15_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_15_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_16 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_16_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_16_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_16_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_17 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_17_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_17_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_17_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_18 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_18_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_18_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_18_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_19 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_19_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_19_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_19_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_20 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_20_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_20_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_20_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_21 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_21_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_21_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_21_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_22 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_22_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_22_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_22_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_23 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_23_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_23_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_23_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_24 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_24_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_24_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_24_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_25 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_25_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_25_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_25_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_26 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_26_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_26_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_26_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_27 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_27_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_27_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_27_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_28 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_28_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_28_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_28_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_29 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_29_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_29_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_29_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_30 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_30_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_30_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_30_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_31 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_31_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_31_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_31_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd128),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a0_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_128_4096_1_4096_128_1_gen
      weight_mem_banks_bank_a1_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_PECoreRun PECore_PECoreRun_inst (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_a(Datapath_for_4_ProductSum_for_acc_5_cmp_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_c(Datapath_for_4_ProductSum_for_acc_5_cmp_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_z(Datapath_for_4_ProductSum_for_acc_5_cmp_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_a(Datapath_for_4_ProductSum_for_acc_5_cmp_1_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_c(Datapath_for_4_ProductSum_for_acc_5_cmp_1_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_z(Datapath_for_4_ProductSum_for_acc_5_cmp_1_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_a(Datapath_for_4_ProductSum_for_acc_5_cmp_2_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_c(Datapath_for_4_ProductSum_for_acc_5_cmp_2_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_z(Datapath_for_4_ProductSum_for_acc_5_cmp_2_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_a(Datapath_for_4_ProductSum_for_acc_5_cmp_3_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_c(Datapath_for_4_ProductSum_for_acc_5_cmp_3_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_z(Datapath_for_4_ProductSum_for_acc_5_cmp_3_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_4_a(Datapath_for_4_ProductSum_for_acc_5_cmp_4_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_4_c(Datapath_for_4_ProductSum_for_acc_5_cmp_4_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_4_z(Datapath_for_4_ProductSum_for_acc_5_cmp_4_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_a(Datapath_for_4_ProductSum_for_acc_5_cmp_5_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_c(Datapath_for_4_ProductSum_for_acc_5_cmp_5_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_en(Datapath_for_4_ProductSum_for_acc_5_cmp_5_en),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_z(Datapath_for_4_ProductSum_for_acc_5_cmp_5_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_6_a(Datapath_for_4_ProductSum_for_acc_5_cmp_6_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_6_c(Datapath_for_4_ProductSum_for_acc_5_cmp_6_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_6_z(Datapath_for_4_ProductSum_for_acc_5_cmp_6_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_7_a(Datapath_for_4_ProductSum_for_acc_5_cmp_7_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_7_c(Datapath_for_4_ProductSum_for_acc_5_cmp_7_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_7_z(Datapath_for_4_ProductSum_for_acc_5_cmp_7_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_8_a(Datapath_for_4_ProductSum_for_acc_5_cmp_8_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_8_c(Datapath_for_4_ProductSum_for_acc_5_cmp_8_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_8_z(Datapath_for_4_ProductSum_for_acc_5_cmp_8_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_9_a(Datapath_for_4_ProductSum_for_acc_5_cmp_9_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_9_c(Datapath_for_4_ProductSum_for_acc_5_cmp_9_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_9_z(Datapath_for_4_ProductSum_for_acc_5_cmp_9_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_10_a(Datapath_for_4_ProductSum_for_acc_5_cmp_10_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_10_c(Datapath_for_4_ProductSum_for_acc_5_cmp_10_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_10_z(Datapath_for_4_ProductSum_for_acc_5_cmp_10_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_11_a(Datapath_for_4_ProductSum_for_acc_5_cmp_11_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_11_c(Datapath_for_4_ProductSum_for_acc_5_cmp_11_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_11_z(Datapath_for_4_ProductSum_for_acc_5_cmp_11_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_12_a(Datapath_for_4_ProductSum_for_acc_5_cmp_12_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_12_c(Datapath_for_4_ProductSum_for_acc_5_cmp_12_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_12_z(Datapath_for_4_ProductSum_for_acc_5_cmp_12_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_13_a(Datapath_for_4_ProductSum_for_acc_5_cmp_13_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_13_c(Datapath_for_4_ProductSum_for_acc_5_cmp_13_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_13_z(Datapath_for_4_ProductSum_for_acc_5_cmp_13_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_14_a(Datapath_for_4_ProductSum_for_acc_5_cmp_14_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_14_c(Datapath_for_4_ProductSum_for_acc_5_cmp_14_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_14_z(Datapath_for_4_ProductSum_for_acc_5_cmp_14_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_15_a(Datapath_for_4_ProductSum_for_acc_5_cmp_15_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_15_c(Datapath_for_4_ProductSum_for_acc_5_cmp_15_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_15_z(Datapath_for_4_ProductSum_for_acc_5_cmp_15_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_16_a(Datapath_for_4_ProductSum_for_acc_5_cmp_16_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_16_c(Datapath_for_4_ProductSum_for_acc_5_cmp_16_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_16_z(Datapath_for_4_ProductSum_for_acc_5_cmp_16_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_17_a(Datapath_for_4_ProductSum_for_acc_5_cmp_17_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_17_c(Datapath_for_4_ProductSum_for_acc_5_cmp_17_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_17_z(Datapath_for_4_ProductSum_for_acc_5_cmp_17_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_18_a(Datapath_for_4_ProductSum_for_acc_5_cmp_18_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_18_c(Datapath_for_4_ProductSum_for_acc_5_cmp_18_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_18_z(Datapath_for_4_ProductSum_for_acc_5_cmp_18_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_19_a(Datapath_for_4_ProductSum_for_acc_5_cmp_19_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_19_c(Datapath_for_4_ProductSum_for_acc_5_cmp_19_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_19_z(Datapath_for_4_ProductSum_for_acc_5_cmp_19_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_20_a(Datapath_for_4_ProductSum_for_acc_5_cmp_20_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_20_c(Datapath_for_4_ProductSum_for_acc_5_cmp_20_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_20_z(Datapath_for_4_ProductSum_for_acc_5_cmp_20_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_a(Datapath_for_4_ProductSum_for_acc_5_cmp_21_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_c(Datapath_for_4_ProductSum_for_acc_5_cmp_21_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_z(Datapath_for_4_ProductSum_for_acc_5_cmp_21_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_22_a(Datapath_for_4_ProductSum_for_acc_5_cmp_22_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_22_c(Datapath_for_4_ProductSum_for_acc_5_cmp_22_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_22_z(Datapath_for_4_ProductSum_for_acc_5_cmp_22_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_23_a(Datapath_for_4_ProductSum_for_acc_5_cmp_23_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_23_c(Datapath_for_4_ProductSum_for_acc_5_cmp_23_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_23_z(Datapath_for_4_ProductSum_for_acc_5_cmp_23_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_24_a(Datapath_for_4_ProductSum_for_acc_5_cmp_24_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_24_c(Datapath_for_4_ProductSum_for_acc_5_cmp_24_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_24_z(Datapath_for_4_ProductSum_for_acc_5_cmp_24_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_25_a(Datapath_for_4_ProductSum_for_acc_5_cmp_25_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_25_c(Datapath_for_4_ProductSum_for_acc_5_cmp_25_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_25_z(Datapath_for_4_ProductSum_for_acc_5_cmp_25_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_26_a(Datapath_for_4_ProductSum_for_acc_5_cmp_26_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_26_c(Datapath_for_4_ProductSum_for_acc_5_cmp_26_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_26_z(Datapath_for_4_ProductSum_for_acc_5_cmp_26_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_27_a(Datapath_for_4_ProductSum_for_acc_5_cmp_27_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_27_c(Datapath_for_4_ProductSum_for_acc_5_cmp_27_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_27_z(Datapath_for_4_ProductSum_for_acc_5_cmp_27_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_28_a(Datapath_for_4_ProductSum_for_acc_5_cmp_28_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_28_c(Datapath_for_4_ProductSum_for_acc_5_cmp_28_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_28_z(Datapath_for_4_ProductSum_for_acc_5_cmp_28_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_29_a(Datapath_for_4_ProductSum_for_acc_5_cmp_29_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_29_c(Datapath_for_4_ProductSum_for_acc_5_cmp_29_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_29_z(Datapath_for_4_ProductSum_for_acc_5_cmp_29_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_30_a(Datapath_for_4_ProductSum_for_acc_5_cmp_30_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_30_c(Datapath_for_4_ProductSum_for_acc_5_cmp_30_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_30_z(Datapath_for_4_ProductSum_for_acc_5_cmp_30_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_31_a(Datapath_for_4_ProductSum_for_acc_5_cmp_31_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_31_c(Datapath_for_4_ProductSum_for_acc_5_cmp_31_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_31_z(Datapath_for_4_ProductSum_for_acc_5_cmp_31_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_5_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_5_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_6_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_6_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_7_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_7_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_8_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_8_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff)
    );
endmodule



