
//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 05:40:36 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [312:0] this_dat;
  output [255:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [255:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_dat[255:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_dat[279:256];
  wire  nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_dat[312];
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd256)) data_data_rsci (
      .d(nl_data_data_rsci_d[255:0]),
      .z(data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d),
      .z(data_rw_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd154),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [312:0] this_dat;
  output [255:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 05:40:31 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [265:0] this_dat;
  output [255:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [255:0] nl_data_data_data_rsci_d;
  assign nl_data_data_data_rsci_d = this_dat[255:0];
  wire [7:0] nl_data_logical_addr_rsci_d;
  assign nl_data_logical_addr_rsci_d = this_dat[265:258];
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd7),
  .width(32'sd256)) data_data_data_rsci (
      .d(nl_data_data_data_rsci_d[255:0]),
      .z(data_data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd9),
  .width(32'sd8)) data_logical_addr_rsci (
      .d(nl_data_logical_addr_rsci_d[7:0]),
      .z(data_logical_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd11),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd153),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [265:0] this_dat;
  output [255:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_data_rsc_z(data_data_data_rsc_z),
      .data_logical_addr_rsc_z(data_logical_addr_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 04:38:53 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [255:0] this_dat;
  reg [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [255:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd13),
  .width(32'sd256)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd152),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd156)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 01:32:50 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd15),
  .width(32'sd1)) data_rsci (
      .d(this_dat),
      .z(data_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd17),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd151),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 05:40:34 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [255:0] this_dat;
  reg [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [255:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd18),
  .width(32'sd256)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd150),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd155)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module PECore_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // spyglass disable SYNTH_5121,W240
    input                s_rst;  // spyglass disable SYNTH_5121,W240
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a; //spyglass disable FlopEConst
                b_reg[0] <= b; //spyglass disable FlopEConst
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> ./PECore_mgc_muladd1_beh.v 
//muladd1
module PECore_mgc_muladd1(a,b,c,cst,d,z);
  // operation is z = a * (b + d) + c + cst
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_cst = 0;
  parameter signd_cst = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_axb = 1;
  parameter add_c = 1;
  parameter add_d = 1;
  parameter use_const = 1;

  function integer is_square_op;
    input integer alen;
  begin
    if (alen > 1) is_square_op = 0;
    else       is_square_op = 1;
  end endfunction

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_cst-1:0] cst; // spyglass disable SYNTH_5121,W240
  input  [width_d-1:0] d;
  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa;
  reg [width_b-signd_b:0] bb;
  reg [width_c-signd_c:0] cc;
  reg [width_d-signd_d:0] dd;
  reg [width_cst-signd_cst:0] cstin;

  localparam width_bd = (width_d) ? 1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b
                                                                          : width_d - signd_d)
                                  : width_b - signd_b;
  localparam is_square = is_square_op(width_a);
  localparam axb_len = (is_square)?width_bd+1+width_bd+1:width_a-signd_a+1+width_bd+1;

  reg [width_bd:0] bd;
  reg [axb_len-1:0] axb;



  // make all inputs signed
  always @(*) aa = signd_a ? a : {1'b0, a};
  always @(*) bb = signd_b ? b : {1'b0, b};
  generate if (width_c != 0) begin
    always @(*) cc = signd_c ? c : {1'b0, c};
  end endgenerate

  generate if (width_d) begin
    if ( !is_square) begin
      (* keep ="true" *) reg [width_d-signd_d:0] d_keep;
      always @(*) d_keep = signd_d ? d : {1'b0, d};
      always @(*) dd = d_keep;
    end else begin
      always @(*) dd = signd_d ? d : {1'b0, d};
    end
  end endgenerate

  always @(*) cstin = signd_cst ? cst : {1'b0, cst};

  // perform pre-adder
  generate
    if (width_d != 0) begin
      if (add_d) begin always @(*)  bd = $signed(bb) + $signed(dd); end
      else       begin always @(*)  bd = $signed(bb) - $signed(dd); end
    end else     begin always @(*)  bd = $signed(bb); end
  endgenerate

  generate
    if (is_square)
      always @(*) axb = $signed(bd) * $signed(bd);
    else
      always @(*) axb = $signed(aa) * $signed(bd);
  endgenerate

  // perform muladd1
  wire [width_z-1:0]  zz;

  generate
    if (use_const) begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc) + $signed(cstin); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc) + $signed(cstin); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb) + $signed(cstin); end else
      if (!add_axb && !add_c && width_c) begin assign zz = $signed(cstin) - $signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb) + $signed(cstin); end else
                                         begin assign zz = $signed(cstin) - $signed(axb); end
    end  else begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb); end else
      if (!add_axb && !add_c && width_c) begin assign zz = -$signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb); end else
                                         begin assign zz = -$signed(axb); end
    end
  endgenerate

  // adjust output
  assign z = zz;
endmodule // mgc_muladd1

//------> ./PECore_mgc_shift_l_beh_v5.v 
module PECore_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./PECore_mgc_mul2add1_pipe_beh.v 
//muladd1
module PECore_mgc_mul2add1_pipe(a,b,b2,c,d,d2,cst,clk,en,a_rst,s_rst,z);
  parameter gentype = 0;
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_b2 = 0;
  parameter signd_b2 = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_d2 = 0;
  parameter signd_d2 = 0;
  parameter width_e = 0;
  parameter signd_e = 0;
  parameter width_z = 0;
  parameter isadd = 1;
  parameter add_b2 = 1;
  parameter add_d2 = 1;
  parameter use_const = 1;
  parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
  parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
  parameter    a_rst_active =  1'b1;  // unused
  parameter    s_rst_active =  1'b1;  // unused
  parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
  parameter integer n_inreg = 32'd0;  // number of input registers

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_b2-1:0] b2; // spyglass disable SYNTH_5121,W240
  input  [width_c-1:0] c;
  input  [width_d-1:0] d;
  input  [width_d2-1:0] d2; // spyglass disable SYNTH_5121,W240
  input  [width_e-1:0] cst; // spyglass disable SYNTH_5121,W240

  input                clk;    // clock
  input                en;     // enable
  input                a_rst;  // spyglass disable SYNTH_5121,W240
  input                s_rst;  // spyglass disable SYNTH_5121,W240

  output [width_z-1:0] z;

  function integer MIN;
    input integer a, b;
  begin
    if (a > b) MIN = b;
    else       MIN = a;
  end endfunction

  function integer f_axb_stages;
    input integer gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d;
  begin
    if (gentype%2==0) begin
      if ((n_inreg > 1) && (width_a>18 | width_b>=19+signd_b | width_c>18 | width_d>=19+signd_d ))
        f_axb_stages = 1;
      else
        f_axb_stages = 0;
    end else begin
      if (n_inreg>1)
        f_axb_stages = 1;
      else
        f_axb_stages = 0;
    end
  end endfunction

  function integer f_cxd_stages;
    input integer gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d;
  begin
    if (gentype%2==0) begin
      f_cxd_stages = 0;
    end else begin
      if (n_inreg>1)
        f_cxd_stages = MIN(n_inreg-1,3);
      else
        f_cxd_stages = 0;
    end
  end endfunction

  function integer f_preadd_stages;
    input integer gentype,n_inreg,width_preaddin;
  begin
    if (gentype%2==0) begin
      f_preadd_stages = 0;
    end else begin
      if (n_inreg>1) begin
        if (width_preaddin>0)
          f_preadd_stages = 1;
        else
          f_preadd_stages = 0;
      end else
        f_preadd_stages = 0;
    end
  end endfunction

  function integer MAX;
    input integer LEFT, RIGHT;
  begin
    if (LEFT > RIGHT) MAX = LEFT;
    else              MAX = RIGHT;
  end endfunction

  function integer PREADDLEN;
    input integer b_len, d_len, width_d;
  begin
    if(width_d>0) PREADDLEN = MAX(b_len,d_len) + 1;
    else        PREADDLEN = b_len;
  end endfunction
  function integer PREADDMULLEN;
    input integer a_len, b_len, d_len, width_d;
  begin
    PREADDMULLEN = a_len + PREADDLEN(b_len,d_len,width_d);
  end endfunction

  localparam axb_stages = f_axb_stages(gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d);
  localparam cxd_stages = f_cxd_stages(gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d);
  localparam preadd_ab_stages = f_preadd_stages(gentype, n_inreg - axb_stages,width_b2);
  localparam preadd_cd_stages = f_preadd_stages(gentype, n_inreg - cxd_stages,width_d2);
  localparam e_stages  = (use_const>1)?n_inreg:0;
  localparam a_stages  = n_inreg - axb_stages;
  localparam b_stages  = n_inreg - axb_stages - preadd_ab_stages;
  localparam c_stages  = n_inreg - cxd_stages;
  localparam d_stages  = n_inreg - cxd_stages - preadd_cd_stages;
  localparam b2_stages  = (width_b2>0)?b_stages:0;
  localparam d2_stages  = (width_d2>0)?d_stages:0;

  localparam a_len    = width_a-signd_a+1;
  localparam b_len    = width_b-signd_b+1;
  localparam b2_len   = width_b2-signd_b2+1;
  localparam c_len    = width_c-signd_c+1;
  localparam d_len    = width_d-signd_d+1;
  localparam d2_len   = width_d2-signd_d2+1;
  localparam e_len    = width_e-signd_e+1;
  localparam bb2_len  = PREADDLEN(b_len, b2_len, width_b2);
  localparam dd2_len  = PREADDLEN(d_len, d2_len, width_d2);
  localparam axb_len  = PREADDMULLEN(a_len, b_len, b2_len, width_b2);
  localparam cxd_len  = PREADDMULLEN(c_len, d_len, d2_len, width_d2);
  localparam z_len    = width_z;

  reg [a_len-1:0]  aa  [a_stages:0];
  reg [b_len-1:0]  bb  [b_stages:0];
  reg [b2_len-1:0] bb2 [b2_stages:0];
  reg [c_len-1:0]  cc  [c_stages:0];
  reg [d_len-1:0]  dd  [d_stages:0];
  reg [d2_len-1:0] dd2 [d2_stages:0];
  reg [e_len-1:0]  ee  [e_stages:0];



  genvar i;

  // make all inputs signed
  always @(*) aa[a_stages] = signd_a ? a : {1'b0, a}; //spyglass disable W164a W164b
  always @(*) bb[b_stages] = signd_b ? b : {1'b0, b}; //spyglass disable W164a W164b
  generate if (width_b2>0) begin
    (* keep ="true" *) reg [b2_len-1:0] b2_keep;
    always @(*) b2_keep = signd_b2 ? b2 : {1'b0, b2}; //spyglass disable W164a W164b
    always @(*) bb2[b2_stages] = b2_keep;
  end endgenerate
  always @(*) cc[c_stages] = signd_c ? c : {1'b0, c}; //spyglass disable W164a W164b
  always @(*) dd[d_stages] = signd_d ? d : {1'b0, d}; //spyglass disable W164a W164b
  generate if (width_d2>0) begin
    (* keep ="true" *) reg [d2_len-1:0] d2_keep;
    always @(*) d2_keep = signd_d2 ? d2 : {1'b0, d2}; //spyglass disable W164a W164b
    always @(*) dd2[d2_stages] = d2_keep;
  end endgenerate

  generate if (use_const>0) begin
    always @(*) ee[e_stages] = signd_e ? cst : {1'b0, cst}; //spyglass disable W164a W164b

    // input registers
    if (e_stages>0) begin
    for(i = e_stages-1; i >= 0; i=i-1) begin:in_pipe_e
      if (clock_edge == 1'b1) begin:pos
        always @(posedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
      end else begin:neg
        always @(negedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
      end
    end end
  end endgenerate
  generate if (a_stages>0) begin
  for(i = a_stages-1; i >= 0; i=i-1) begin:in_pipe_a
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (b_stages>0) begin
  for(i = b_stages-1; i >= 0; i=i-1) begin:in_pipe_b
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];
    end
  end end endgenerate
  generate if (c_stages>0) begin
  for(i = c_stages-1; i >= 0; i=i-1) begin:in_pipe_c
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (d_stages>0) begin
  for(i = d_stages-1; i >= 0; i=i-1) begin:in_pipe_d
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) dd[i] <= dd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) dd[i] <= dd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (b2_stages>0) begin
  for(i = b2_stages-1; i >= 0; i=i-1) begin:in_pipe_b2
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb2[i] <= bb2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb2[i] <= bb2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (d2_stages>0) begin
  for(i = d2_stages-1; i >= 0; i=i-1) begin:in_pipe_d2
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) dd2[i] <= dd2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) dd2[i] <= dd2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg [bb2_len-1:0] b_bb2[preadd_ab_stages:0];
  reg [dd2_len-1:0] d_dd2[preadd_cd_stages:0];

  //perform first preadd
  generate
    if (width_b2>0) begin
      if (add_b2) begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]) + $signed(bb2[0]); end
      else        begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]) - $signed(bb2[0]); end
    end else      begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]); end
  endgenerate
  generate if (preadd_ab_stages>0) begin
  for(i = preadd_ab_stages-1; i >= 0; i=i-1) begin:preaddab_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) b_bb2[i] <= b_bb2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) b_bb2[i] <= b_bb2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  //perform second preadd
  generate
    if (width_d2>0) begin
      if (add_d2) begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]) + $signed(dd2[0]); end
      else        begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]) - $signed(dd2[0]); end
    end else      begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]); end
  endgenerate
  generate if (preadd_cd_stages>0) begin
  for(i = preadd_cd_stages-1; i >= 0; i=i-1) begin:preaddcd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) d_dd2[i] <= d_dd2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) d_dd2[i] <= d_dd2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // perform first multiplication
  reg [axb_len-1:0] axb[axb_stages:0];

  always @(*) axb[axb_stages] = $signed(aa[0]) * $signed(b_bb2[0]);
  generate if (axb_stages>0) begin
  for(i = axb_stages-1; i >= 0; i=i-1) begin:axb_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];
    end
  end end endgenerate

  // perform second multiplication
  reg [cxd_len-1:0] cxd[cxd_stages:0];

  always @(*) cxd[cxd_stages] = $signed(cc[0]) * $signed(d_dd2[0]);
  generate if (cxd_stages>0) begin
  for(i = cxd_stages-1; i >= 0; i=i-1) begin:cxd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cxd[i] <= cxd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cxd[i] <= cxd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg [z_len-1:0]  zz[stages-1:0];
  generate
    if (use_const>1) begin
      reg [z_len-1:0] aux_val;
      if ( isadd) begin
        always @(*) aux_val = $signed(axb[0]) + $signed(cxd[0]);
      end else begin
        always @(*) aux_val = $signed(axb[0]) - $signed(cxd[0]);
      end
      always @(*) zz[stages-1] = $signed(ee[0]) + $signed(aux_val) ;
    end else begin
      if (use_const>0) begin
        if ( isadd) begin always @(*) zz[stages-1] = $signed(axb[0]) + $signed(cxd[0]) + $signed(ee[0]); end else
                    begin always @(*) zz[stages-1] = $signed(axb[0]) - $signed(cxd[0]) + $signed(ee[0]); end
      end else begin
        if ( isadd) begin always @(*) zz[stages-1] = $signed(axb[0]) + $signed(cxd[0]); end else
                    begin always @(*) zz[stages-1] = $signed(axb[0]) - $signed(cxd[0]); end
      end
    end
  endgenerate

  // Output registers:
  generate if (stages>1) begin
  for(i = stages-2; i >= 0; i=i-1) begin:out_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // adjust output
  assign z = zz[0];
endmodule // mgc_mul2add1_pipe

//------> /cad/mentor/2024.2_1/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)
// suppress_sim_read_addr_range_errs:  0 - report errors  1 - suppress errors

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 ,
  parameter suppress_sim_read_addr_range_errs = 1 
  
)( clk,clken,d,q,radr,re,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input  re;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" , syn_ramstyle = "block" *)
  reg [data_width-1:0] mem [depth-1:0];
  integer j;
  initial for (j = 0; j < depth; j = j + 1) mem[j] = 0;
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr READ_ENABLE re
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg re_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
          re_reg <= re;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./PECore.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 05:54:34 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_256_4096_1_4096_256_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_256_4096_1_4096_256_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [255:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [255:0] d;
  output [11:0] wadr;
  input clken_d;
  input [255:0] d_d;
  output [255:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_256_4096_1_4096_256_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_256_4096_1_4096_256_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [255:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [255:0] d;
  output [11:0] wadr;
  input clken_d;
  input [255:0] d_d;
  output [255:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_256_4096_1_4096_256_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_256_4096_1_4096_256_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [255:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [255:0] d;
  output [11:0] wadr;
  input clken_d;
  input [255:0] d_d;
  output [255:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_256_4096_1_4096_256_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_256_4096_1_4096_256_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [255:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [255:0] d;
  output [11:0] wadr;
  input clken_d;
  input [255:0] d_d;
  output [255:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_256_4096_1_4096_256_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_256_4096_1_4096_256_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [255:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [255:0] d;
  output [11:0] wadr;
  input clken_d;
  input [255:0] d_d;
  output [255:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_256_4096_1_4096_256_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_256_4096_1_4096_256_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [255:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [255:0] d;
  output [11:0] wadr;
  input clken_d;
  input [255:0] d_d;
  output [255:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_256_4096_1_4096_256_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_256_4096_1_4096_256_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [255:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [255:0] d;
  output [11:0] wadr;
  input clken_d;
  input [255:0] d_d;
  output [255:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_256_4096_1_4096_256_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_256_4096_1_4096_256_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [255:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [255:0] d;
  output [11:0] wadr;
  input clken_d;
  input [255:0] d_d;
  output [255:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_PECoreRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_PECoreRun_fsm (
  clk, rst, PECoreRun_wen, fsm_output
);
  input clk;
  input rst;
  input PECoreRun_wen;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for PECore_PECore_PECoreRun_PECoreRun_fsm_1
  parameter
    PECoreRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : PECore_PECore_PECoreRun_PECoreRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // PECoreRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= PECoreRun_rlp_C_0;
    end
    else if ( PECoreRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_staller
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_staller (
  clk, rst, PECoreRun_wen, PECoreRun_wten, act_port_Push_mioi_wen_comp, rva_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PECoreRun_wen;
  output PECoreRun_wten;
  input act_port_Push_mioi_wen_comp;
  input rva_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg PECoreRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign PECoreRun_wen = act_port_Push_mioi_wen_comp & rva_out_Push_mioi_wen_comp;
  assign PECoreRun_wten = PECoreRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECoreRun_wten_reg <= 1'b0;
    end
    else begin
      PECoreRun_wten_reg <= ~ PECoreRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_wait_dp (
  weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      Datapath_for_4_ProductSum_for_acc_9_cmp_en, Datapath_for_4_ProductSum_for_acc_9_cmp_1_en,
      PECoreRun_wen, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg,
      PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo, PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg,
      PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en, PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_1,
      PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg_1, PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en,
      Datapath_for_4_ProductSum_for_acc_9_cmp_cgo, Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg,
      Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_1, Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg_1
);
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output Datapath_for_4_ProductSum_for_acc_9_cmp_en;
  output Datapath_for_4_ProductSum_for_acc_9_cmp_1_en;
  input PECoreRun_wen;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg;
  input PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo;
  input PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg;
  output PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en;
  input PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_1;
  input PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg_1;
  output PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en;
  input Datapath_for_4_ProductSum_for_acc_9_cmp_cgo;
  input Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg;
  input Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_1;
  input Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg_1;



  // Interconnect Declarations for Component Instantiations 
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg);
  assign PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en = PECoreRun_wen & (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo
      | PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg);
  assign PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en = PECoreRun_wen & (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_1
      | PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg_1);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_en = ~(PECoreRun_wen & (Datapath_for_4_ProductSum_for_acc_9_cmp_cgo
      | Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg));
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_en = ~(PECoreRun_wen & (Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_1
      | Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg_1));
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  PECoreRun_wen, rva_out_Push_mioi_oswt, rva_out_Push_mioi_biwt, rva_out_Push_mioi_bdwt,
      rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & PECoreRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt)
      & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & rva_out_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt,
      start_PopNB_mioi_biwt_pff, start_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_biwt_pff;
  input start_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & PECoreRun_wen;
  assign start_PopNB_mioi_biwt = (~ PECoreRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_biwt_pff = PECoreRun_wen & start_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp (
  clk, rst, act_port_Push_mioi_oswt, act_port_Push_mioi_wen_comp, act_port_Push_mioi_biwt,
      act_port_Push_mioi_bdwt, act_port_Push_mioi_bcwt
);
  input clk;
  input rst;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input act_port_Push_mioi_biwt;
  input act_port_Push_mioi_bdwt;
  output act_port_Push_mioi_bcwt;
  reg act_port_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_wen_comp = (~ act_port_Push_mioi_oswt) | act_port_Push_mioi_biwt
      | act_port_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_Push_mioi_bcwt <= ~((~(act_port_Push_mioi_bcwt | act_port_Push_mioi_biwt))
          | act_port_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl (
  PECoreRun_wen, act_port_Push_mioi_oswt, act_port_Push_mioi_biwt, act_port_Push_mioi_bdwt,
      act_port_Push_mioi_bcwt, act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      act_port_Push_mioi_ccs_ccore_done_sync_vld, act_port_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_biwt;
  output act_port_Push_mioi_bdwt;
  input act_port_Push_mioi_bcwt;
  output act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input act_port_Push_mioi_ccs_ccore_done_sync_vld;
  input act_port_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_bdwt = act_port_Push_mioi_oswt & PECoreRun_wen;
  assign act_port_Push_mioi_biwt = act_port_Push_mioi_oswt & (~ act_port_Push_mioi_bcwt)
      & act_port_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & act_port_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
    (
  clk, rst, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt,
      input_port_PopNB_mioi_return_rsc_z_mxwt, input_port_PopNB_mioi_biwt, input_port_PopNB_mioi_bdwt,
      input_port_PopNB_mioi_data_data_data_rsc_z, input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [255:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_biwt;
  input input_port_PopNB_mioi_bdwt;
  input [255:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  input [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  input input_port_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg input_port_PopNB_mioi_bcwt;
  reg [255:0] input_port_PopNB_mioi_data_data_data_rsc_z_bfwt;
  reg [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt;
  reg input_port_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_data_data_data_rsc_z_mxwt = MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z,
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt = MUX_v_8_2_2(input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z,
      input_port_PopNB_mioi_return_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      input_port_PopNB_mioi_bcwt <= ~((~(input_port_PopNB_mioi_bcwt | input_port_PopNB_mioi_biwt))
          | input_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= 8'b00000000;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( input_port_PopNB_mioi_biwt ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= input_port_PopNB_mioi_data_data_data_rsc_z;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= input_port_PopNB_mioi_data_logical_addr_rsc_z;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= input_port_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input  sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
    (
  PECoreRun_wen, PECoreRun_wten, input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_biwt,
      input_port_PopNB_mioi_bdwt, input_port_PopNB_mioi_biwt_pff, input_port_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output input_port_PopNB_mioi_biwt;
  output input_port_PopNB_mioi_bdwt;
  output input_port_PopNB_mioi_biwt_pff;
  input input_port_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_bdwt = input_port_PopNB_mioi_oswt & PECoreRun_wen;
  assign input_port_PopNB_mioi_biwt = (~ PECoreRun_wten) & input_port_PopNB_mioi_oswt;
  assign input_port_PopNB_mioi_biwt_pff = PECoreRun_wen & input_port_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [255:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [255:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [255:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  reg [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_256_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_20_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4, rva_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= 20'b00000000000000000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input  sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & PECoreRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ PECoreRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = PECoreRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, PECoreRun_wen, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_PECoreRun, rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [255:0] rva_out_dat;
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [255:0] rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_oswt_pff(rva_out_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi (
  clk, rst, start_vld, start_rdy, start_dat, PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_vld(start_vld),
      .this_rdy(start_rdy),
      .this_dat(start_dat),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_biwt_pff(start_PopNB_mioi_biwt_iff),
      .start_PopNB_mioi_oswt_pff(start_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi (
  clk, rst, act_port_vld, act_port_rdy, act_port_dat, PECoreRun_wen, act_port_Push_mioi_oswt,
      act_port_Push_mioi_wen_comp, act_port_Push_mioi_m_data_rsc_dat_PECoreRun, act_port_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input [255:0] act_port_Push_mioi_m_data_rsc_dat_PECoreRun;
  input act_port_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_port_Push_mioi_biwt;
  wire act_port_Push_mioi_bdwt;
  wire act_port_Push_mioi_bcwt;
  wire act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire act_port_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push  act_port_Push_mioi
      (
      .this_vld(act_port_vld),
      .this_rdy(act_port_rdy),
      .this_dat(act_port_dat),
      .m_data_rsc_dat(act_port_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt),
      .act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .act_port_Push_mioi_ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .act_port_Push_mioi_oswt_pff(act_port_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi (
  clk, rst, input_port_vld, input_port_rdy, input_port_dat, PECoreRun_wen, PECoreRun_wten,
      input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt, input_port_PopNB_mioi_return_rsc_z_mxwt,
      input_port_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input input_port_vld;
  output input_port_rdy;
  input [265:0] input_port_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output [255:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_port_PopNB_mioi_biwt;
  wire input_port_PopNB_mioi_bdwt;
  wire [255:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  wire input_port_PopNB_mioi_return_rsc_z;
  wire input_port_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB  input_port_PopNB_mioi
      (
      .this_vld(input_port_vld),
      .this_rdy(input_port_rdy),
      .this_dat(input_port_dat),
      .data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .return_rsc_z(input_port_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(input_port_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(input_port_PopNB_mioi_oswt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_biwt_pff(input_port_PopNB_mioi_biwt_iff),
      .input_port_PopNB_mioi_oswt_pff(input_port_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .input_port_PopNB_mioi_return_rsc_z(input_port_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt,
      rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [312:0] rva_in_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [255:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [255:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG, weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d, Datapath_for_4_ProductSum_for_acc_9_cmp_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_c, Datapath_for_4_ProductSum_for_acc_9_cmp_en,
      Datapath_for_4_ProductSum_for_acc_9_cmp_z, Datapath_for_4_ProductSum_for_acc_9_cmp_1_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_1_b, Datapath_for_4_ProductSum_for_acc_9_cmp_1_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_1_d, Datapath_for_4_ProductSum_for_acc_9_cmp_1_en,
      Datapath_for_4_ProductSum_for_acc_9_cmp_1_z, Datapath_for_4_ProductSum_for_acc_9_cmp_2_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_2_b, Datapath_for_4_ProductSum_for_acc_9_cmp_2_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_2_d, Datapath_for_4_ProductSum_for_acc_9_cmp_2_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_3_a, Datapath_for_4_ProductSum_for_acc_9_cmp_3_b,
      Datapath_for_4_ProductSum_for_acc_9_cmp_3_c, Datapath_for_4_ProductSum_for_acc_9_cmp_3_d,
      Datapath_for_4_ProductSum_for_acc_9_cmp_3_z, Datapath_for_4_ProductSum_for_acc_9_cmp_4_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_4_b, Datapath_for_4_ProductSum_for_acc_9_cmp_4_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_4_d, Datapath_for_4_ProductSum_for_acc_9_cmp_4_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_5_a, Datapath_for_4_ProductSum_for_acc_9_cmp_5_b,
      Datapath_for_4_ProductSum_for_acc_9_cmp_5_c, Datapath_for_4_ProductSum_for_acc_9_cmp_5_d,
      Datapath_for_4_ProductSum_for_acc_9_cmp_5_z, Datapath_for_4_ProductSum_for_acc_9_cmp_6_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_6_b, Datapath_for_4_ProductSum_for_acc_9_cmp_6_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_6_d, Datapath_for_4_ProductSum_for_acc_9_cmp_6_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_7_a, Datapath_for_4_ProductSum_for_acc_9_cmp_7_b,
      Datapath_for_4_ProductSum_for_acc_9_cmp_7_c, Datapath_for_4_ProductSum_for_acc_9_cmp_7_d,
      Datapath_for_4_ProductSum_for_acc_9_cmp_7_z, Datapath_for_4_ProductSum_for_acc_9_cmp_8_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_8_c, Datapath_for_4_ProductSum_for_acc_9_cmp_8_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_9_a, Datapath_for_4_ProductSum_for_acc_9_cmp_9_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_9_z, Datapath_for_4_ProductSum_for_acc_9_cmp_10_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_10_c, Datapath_for_4_ProductSum_for_acc_9_cmp_10_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_11_a, Datapath_for_4_ProductSum_for_acc_9_cmp_11_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_11_z, Datapath_for_4_ProductSum_for_acc_9_cmp_12_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_12_c, Datapath_for_4_ProductSum_for_acc_9_cmp_12_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_13_a, Datapath_for_4_ProductSum_for_acc_9_cmp_13_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_13_z, Datapath_for_4_ProductSum_for_acc_9_cmp_14_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_14_c, Datapath_for_4_ProductSum_for_acc_9_cmp_14_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_15_a, Datapath_for_4_ProductSum_for_acc_9_cmp_15_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_15_z, Datapath_for_4_ProductSum_for_acc_9_cmp_16_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_16_c, Datapath_for_4_ProductSum_for_acc_9_cmp_16_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_17_a, Datapath_for_4_ProductSum_for_acc_9_cmp_17_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_17_z, Datapath_for_4_ProductSum_for_acc_9_cmp_18_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_18_c, Datapath_for_4_ProductSum_for_acc_9_cmp_18_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_19_a, Datapath_for_4_ProductSum_for_acc_9_cmp_19_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_19_z, Datapath_for_4_ProductSum_for_acc_9_cmp_20_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_20_c, Datapath_for_4_ProductSum_for_acc_9_cmp_20_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_21_a, Datapath_for_4_ProductSum_for_acc_9_cmp_21_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_21_z, Datapath_for_4_ProductSum_for_acc_9_cmp_22_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_22_c, Datapath_for_4_ProductSum_for_acc_9_cmp_22_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_23_a, Datapath_for_4_ProductSum_for_acc_9_cmp_23_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_23_z, Datapath_for_4_ProductSum_for_acc_9_cmp_24_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_24_c, Datapath_for_4_ProductSum_for_acc_9_cmp_24_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_25_a, Datapath_for_4_ProductSum_for_acc_9_cmp_25_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_25_z, Datapath_for_4_ProductSum_for_acc_9_cmp_26_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_26_c, Datapath_for_4_ProductSum_for_acc_9_cmp_26_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_27_a, Datapath_for_4_ProductSum_for_acc_9_cmp_27_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_27_z, Datapath_for_4_ProductSum_for_acc_9_cmp_28_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_28_c, Datapath_for_4_ProductSum_for_acc_9_cmp_28_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_29_a, Datapath_for_4_ProductSum_for_acc_9_cmp_29_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_29_z, Datapath_for_4_ProductSum_for_acc_9_cmp_30_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_30_c, Datapath_for_4_ProductSum_for_acc_9_cmp_30_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_31_a, Datapath_for_4_ProductSum_for_acc_9_cmp_31_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_31_z, Datapath_for_4_ProductSum_for_acc_9_cmp_32_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_32_c, Datapath_for_4_ProductSum_for_acc_9_cmp_32_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_33_a, Datapath_for_4_ProductSum_for_acc_9_cmp_33_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_33_z, Datapath_for_4_ProductSum_for_acc_9_cmp_34_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_34_c, Datapath_for_4_ProductSum_for_acc_9_cmp_34_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_35_a, Datapath_for_4_ProductSum_for_acc_9_cmp_35_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_35_z, Datapath_for_4_ProductSum_for_acc_9_cmp_36_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_36_c, Datapath_for_4_ProductSum_for_acc_9_cmp_36_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_37_a, Datapath_for_4_ProductSum_for_acc_9_cmp_37_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_37_z, Datapath_for_4_ProductSum_for_acc_9_cmp_38_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_38_c, Datapath_for_4_ProductSum_for_acc_9_cmp_38_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_39_a, Datapath_for_4_ProductSum_for_acc_9_cmp_39_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_39_z, Datapath_for_4_ProductSum_for_acc_9_cmp_40_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_40_c, Datapath_for_4_ProductSum_for_acc_9_cmp_40_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_41_a, Datapath_for_4_ProductSum_for_acc_9_cmp_41_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_41_z, Datapath_for_4_ProductSum_for_acc_9_cmp_42_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_42_c, Datapath_for_4_ProductSum_for_acc_9_cmp_42_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_43_a, Datapath_for_4_ProductSum_for_acc_9_cmp_43_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_43_z, Datapath_for_4_ProductSum_for_acc_9_cmp_44_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_44_c, Datapath_for_4_ProductSum_for_acc_9_cmp_44_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_45_a, Datapath_for_4_ProductSum_for_acc_9_cmp_45_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_45_z, Datapath_for_4_ProductSum_for_acc_9_cmp_46_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_46_c, Datapath_for_4_ProductSum_for_acc_9_cmp_46_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_47_a, Datapath_for_4_ProductSum_for_acc_9_cmp_47_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_47_z, Datapath_for_4_ProductSum_for_acc_9_cmp_48_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_48_c, Datapath_for_4_ProductSum_for_acc_9_cmp_48_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_49_a, Datapath_for_4_ProductSum_for_acc_9_cmp_49_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_49_z, Datapath_for_4_ProductSum_for_acc_9_cmp_50_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_50_c, Datapath_for_4_ProductSum_for_acc_9_cmp_50_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_51_a, Datapath_for_4_ProductSum_for_acc_9_cmp_51_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_51_z, Datapath_for_4_ProductSum_for_acc_9_cmp_52_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_52_c, Datapath_for_4_ProductSum_for_acc_9_cmp_52_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_53_a, Datapath_for_4_ProductSum_for_acc_9_cmp_53_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_53_z, Datapath_for_4_ProductSum_for_acc_9_cmp_54_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_54_c, Datapath_for_4_ProductSum_for_acc_9_cmp_54_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_55_a, Datapath_for_4_ProductSum_for_acc_9_cmp_55_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_55_z, Datapath_for_4_ProductSum_for_acc_9_cmp_56_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_56_c, Datapath_for_4_ProductSum_for_acc_9_cmp_56_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_57_a, Datapath_for_4_ProductSum_for_acc_9_cmp_57_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_57_z, Datapath_for_4_ProductSum_for_acc_9_cmp_58_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_58_c, Datapath_for_4_ProductSum_for_acc_9_cmp_58_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_59_a, Datapath_for_4_ProductSum_for_acc_9_cmp_59_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_59_z, Datapath_for_4_ProductSum_for_acc_9_cmp_60_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_60_c, Datapath_for_4_ProductSum_for_acc_9_cmp_60_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_61_a, Datapath_for_4_ProductSum_for_acc_9_cmp_61_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_61_z, Datapath_for_4_ProductSum_for_acc_9_cmp_62_a,
      Datapath_for_4_ProductSum_for_acc_9_cmp_62_c, Datapath_for_4_ProductSum_for_acc_9_cmp_62_z,
      Datapath_for_4_ProductSum_for_acc_9_cmp_63_a, Datapath_for_4_ProductSum_for_acc_9_cmp_63_c,
      Datapath_for_4_ProductSum_for_acc_9_cmp_63_z, Datapath_for_4_ProductSum_for_acc_9_cmp_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_pff, Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_pff,
      Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff, weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [265:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [312:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [255:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output [255:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  input [255:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output [255:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  input [255:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output [255:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  input [255:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output [255:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  input [255:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output [255:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  input [255:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output [255:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  input [255:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output [255:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  input [255:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output [255:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  input [255:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_c;
  output Datapath_for_4_ProductSum_for_acc_9_cmp_en;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_b;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_c;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_d;
  output Datapath_for_4_ProductSum_for_acc_9_cmp_1_en;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_b;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_c;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_d;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_b;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_c;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_d;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_b;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_c;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_d;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_b;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_c;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_d;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_b;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_c;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_d;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_b;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_c;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_d;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_a;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_c;
  input [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_z;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_pff;
  output [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff;


  // Interconnect Declarations
  wire PECoreRun_wen;
  wire PECoreRun_wten;
  wire [255:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [255:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  wire input_port_PopNB_mioi_return_rsc_z_mxwt;
  wire act_port_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_z;
  wire PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_z;
  wire [42:0] PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_z;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
  wire fsm_output;
  wire pe_config_UpdateManagerCounter_if_if_unequal_tmp;
  wire [7:0] weight_mem_write_arbxbar_xbar_for_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_5_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp;
  wire while_mux_1477_tmp;
  wire while_mux_1476_tmp;
  wire while_mux_1475_tmp;
  wire while_mux_1474_tmp;
  wire while_mux_1473_tmp;
  wire while_mux_1472_tmp;
  wire while_mux_1471_tmp;
  wire while_mux_1470_tmp;
  wire while_mux_1469_tmp;
  wire while_mux_1468_tmp;
  wire while_mux_1467_tmp;
  wire while_mux_1466_tmp;
  wire while_mux_1465_tmp;
  wire while_mux_1464_tmp;
  wire while_mux_1456_tmp;
  wire while_mux_1454_tmp;
  wire while_mux_1451_tmp;
  wire while_mux_1450_tmp;
  wire while_mux_1445_tmp;
  wire while_mux_1435_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_125_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_30_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp;
  wire weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
  wire while_and_46_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  wire and_dcpl_6;
  wire and_dcpl_7;
  wire and_dcpl_8;
  wire and_dcpl_24;
  wire and_dcpl_40;
  wire or_tmp;
  wire and_dcpl_45;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_76;
  wire and_dcpl_85;
  wire and_dcpl_87;
  wire and_dcpl_89;
  wire and_dcpl_91;
  wire or_dcpl_32;
  wire and_dcpl_93;
  wire and_dcpl_95;
  wire and_dcpl_97;
  wire and_dcpl_99;
  wire and_dcpl_101;
  wire or_dcpl_47;
  wire or_dcpl_48;
  wire or_dcpl_50;
  wire or_dcpl_53;
  wire and_dcpl_123;
  wire and_dcpl_124;
  wire and_dcpl_125;
  wire and_dcpl_126;
  wire and_dcpl_127;
  wire and_dcpl_128;
  wire and_dcpl_129;
  wire and_dcpl_130;
  wire and_dcpl_133;
  wire and_dcpl_137;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire and_dcpl_156;
  wire and_dcpl_157;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire and_dcpl_161;
  wire and_dcpl_162;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_167;
  wire and_dcpl_168;
  wire and_dcpl_169;
  wire and_dcpl_172;
  wire and_dcpl_176;
  wire and_dcpl_179;
  wire and_dcpl_180;
  wire or_dcpl_121;
  wire or_dcpl_126;
  wire or_dcpl_129;
  wire and_dcpl_183;
  wire and_dcpl_186;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire and_dcpl_191;
  wire and_dcpl_195;
  wire or_tmp_35;
  wire and_dcpl_226;
  wire and_dcpl_230;
  wire and_dcpl_231;
  wire and_dcpl_241;
  wire and_dcpl_253;
  wire and_dcpl_258;
  wire not_tmp_139;
  wire mux_tmp_46;
  wire and_dcpl_274;
  wire and_dcpl_282;
  wire and_dcpl_284;
  wire and_dcpl_312;
  wire and_dcpl_313;
  wire and_dcpl_320;
  wire and_dcpl_321;
  wire mux_tmp_51;
  wire or_tmp_59;
  wire and_dcpl_325;
  wire and_dcpl_343;
  wire and_dcpl_344;
  wire and_dcpl_347;
  wire and_dcpl_348;
  wire or_dcpl_177;
  wire or_dcpl_178;
  wire or_dcpl_179;
  wire or_dcpl_180;
  wire or_dcpl_181;
  wire or_dcpl_182;
  wire or_dcpl_185;
  wire or_dcpl_187;
  wire or_dcpl_188;
  wire or_dcpl_189;
  wire or_dcpl_191;
  wire or_dcpl_192;
  wire or_dcpl_193;
  wire or_dcpl_195;
  wire or_dcpl_196;
  wire or_dcpl_197;
  wire or_dcpl_199;
  wire or_dcpl_200;
  wire or_dcpl_201;
  wire or_dcpl_203;
  wire or_dcpl_205;
  wire or_dcpl_207;
  wire or_dcpl_209;
  wire or_dcpl_210;
  wire or_dcpl_211;
  wire or_dcpl_213;
  wire or_dcpl_215;
  wire or_dcpl_217;
  wire or_dcpl_219;
  wire or_dcpl_220;
  wire or_dcpl_221;
  wire or_dcpl_223;
  wire or_dcpl_225;
  wire or_dcpl_227;
  wire or_dcpl_229;
  wire or_dcpl_230;
  wire or_dcpl_232;
  wire or_dcpl_234;
  wire or_dcpl_236;
  wire or_dcpl_238;
  wire or_dcpl_239;
  wire or_dcpl_241;
  wire or_dcpl_243;
  wire or_dcpl_245;
  wire or_dcpl_247;
  wire or_dcpl_248;
  wire or_dcpl_250;
  wire or_dcpl_252;
  wire or_dcpl_254;
  wire or_dcpl_256;
  wire or_dcpl_257;
  wire or_dcpl_259;
  wire or_dcpl_261;
  wire or_dcpl_263;
  wire or_dcpl_265;
  wire or_dcpl_266;
  wire or_dcpl_267;
  wire or_dcpl_269;
  wire or_dcpl_270;
  wire or_dcpl_272;
  wire or_dcpl_273;
  wire or_dcpl_275;
  wire or_dcpl_276;
  wire or_dcpl_278;
  wire or_dcpl_280;
  wire or_dcpl_282;
  wire or_dcpl_284;
  wire or_dcpl_286;
  wire or_dcpl_288;
  wire or_dcpl_290;
  wire or_dcpl_292;
  wire or_dcpl_294;
  wire or_dcpl_296;
  wire or_dcpl_298;
  wire or_dcpl_300;
  wire or_dcpl_302;
  wire or_dcpl_304;
  wire or_dcpl_306;
  wire or_dcpl_308;
  wire or_dcpl_310;
  wire or_dcpl_312;
  wire or_dcpl_314;
  wire or_dcpl_316;
  wire or_dcpl_318;
  wire or_dcpl_320;
  wire or_dcpl_322;
  wire or_dcpl_324;
  wire or_dcpl_326;
  wire or_dcpl_328;
  wire or_dcpl_330;
  wire or_dcpl_332;
  wire or_dcpl_336;
  wire or_dcpl_401;
  wire or_dcpl_402;
  wire or_dcpl_403;
  wire or_dcpl_405;
  wire or_dcpl_406;
  wire or_dcpl_408;
  wire or_dcpl_409;
  wire or_dcpl_411;
  wire or_dcpl_412;
  wire or_dcpl_414;
  wire or_dcpl_416;
  wire or_dcpl_418;
  wire or_dcpl_420;
  wire or_dcpl_422;
  wire or_dcpl_424;
  wire or_dcpl_426;
  wire or_dcpl_428;
  wire or_dcpl_430;
  wire or_dcpl_432;
  wire or_dcpl_434;
  wire or_dcpl_436;
  wire or_dcpl_438;
  wire or_dcpl_440;
  wire or_dcpl_442;
  wire or_dcpl_444;
  wire or_dcpl_446;
  wire or_dcpl_448;
  wire or_dcpl_450;
  wire or_dcpl_452;
  wire or_dcpl_454;
  wire or_dcpl_456;
  wire or_dcpl_458;
  wire or_dcpl_460;
  wire or_dcpl_462;
  wire or_dcpl_464;
  wire or_dcpl_466;
  wire or_dcpl_468;
  wire or_dcpl_470;
  wire or_dcpl_471;
  wire or_dcpl_472;
  wire or_dcpl_474;
  wire or_dcpl_475;
  wire or_dcpl_477;
  wire or_dcpl_478;
  wire or_dcpl_480;
  wire or_dcpl_481;
  wire or_dcpl_483;
  wire or_dcpl_485;
  wire or_dcpl_487;
  wire or_dcpl_489;
  wire or_dcpl_491;
  wire or_dcpl_493;
  wire or_dcpl_495;
  wire or_dcpl_497;
  wire or_dcpl_499;
  wire or_dcpl_501;
  wire or_dcpl_503;
  wire or_dcpl_505;
  wire or_dcpl_507;
  wire or_dcpl_509;
  wire or_dcpl_511;
  wire or_dcpl_513;
  wire or_dcpl_515;
  wire or_dcpl_517;
  wire or_dcpl_519;
  wire or_dcpl_521;
  wire or_dcpl_523;
  wire or_dcpl_525;
  wire or_dcpl_527;
  wire or_dcpl_529;
  wire or_dcpl_531;
  wire or_dcpl_533;
  wire or_dcpl_535;
  wire or_dcpl_537;
  wire and_dcpl_367;
  wire and_dcpl_371;
  wire and_dcpl_372;
  wire and_dcpl_380;
  wire and_dcpl_395;
  wire and_dcpl_408;
  wire and_dcpl_423;
  wire and_dcpl_444;
  wire or_tmp_68;
  wire and_dcpl_457;
  wire or_dcpl_606;
  wire and_dcpl_468;
  wire and_dcpl_488;
  wire and_dcpl_489;
  wire mux_tmp_69;
  wire and_dcpl_495;
  wire and_dcpl_530;
  wire and_dcpl_532;
  wire or_tmp_75;
  wire or_tmp_76;
  wire or_tmp_78;
  wire and_dcpl_544;
  wire and_tmp_2;
  wire and_dcpl_546;
  wire and_tmp_3;
  wire and_tmp_4;
  wire and_tmp_5;
  wire and_tmp_6;
  wire and_tmp_7;
  wire or_tmp_111;
  wire and_tmp_8;
  wire and_tmp_9;
  wire and_dcpl_567;
  wire and_dcpl_568;
  wire or_dcpl_633;
  wire and_dcpl_584;
  wire and_dcpl_588;
  wire and_dcpl_590;
  wire or_dcpl_636;
  wire or_dcpl_637;
  wire or_dcpl_648;
  wire or_dcpl_649;
  wire and_dcpl_621;
  wire and_dcpl_635;
  wire or_dcpl_700;
  wire and_dcpl_657;
  wire and_dcpl_664;
  wire and_dcpl_674;
  wire and_dcpl_675;
  wire or_dcpl_706;
  wire or_tmp_131;
  wire or_tmp_133;
  wire mux_tmp_126;
  wire nor_tmp_45;
  wire or_tmp_135;
  wire or_tmp_136;
  wire or_tmp_137;
  wire or_tmp_139;
  wire nor_tmp_51;
  wire or_tmp_141;
  wire or_tmp_142;
  wire or_tmp_143;
  wire or_tmp_145;
  wire or_tmp_149;
  wire or_tmp_150;
  wire or_tmp_151;
  wire or_tmp_155;
  wire or_tmp_156;
  wire or_tmp_157;
  wire and_dcpl_680;
  wire or_tmp_174;
  wire or_tmp_177;
  wire or_tmp_179;
  wire or_tmp_181;
  wire mux_tmp_149;
  wire mux_tmp_152;
  wire mux_tmp_155;
  wire nor_tmp_83;
  wire or_tmp_186;
  wire or_tmp_191;
  wire or_tmp_194;
  wire mux_tmp_162;
  wire or_tmp_198;
  wire nor_tmp_90;
  wire or_tmp_204;
  wire nor_tmp_93;
  wire or_tmp_210;
  wire and_dcpl_683;
  wire or_tmp_219;
  wire or_tmp_224;
  wire or_dcpl_710;
  wire and_dcpl_685;
  wire or_tmp_226;
  wire or_tmp_228;
  wire and_dcpl_686;
  wire and_dcpl_687;
  wire and_dcpl_688;
  wire and_dcpl_689;
  wire mux_tmp_187;
  wire mux_tmp_188;
  wire mux_tmp_189;
  wire and_dcpl_690;
  wire and_dcpl_696;
  wire nor_tmp_107;
  wire nor_tmp_109;
  wire or_dcpl_711;
  wire nand_tmp_9;
  wire nand_tmp_10;
  wire and_dcpl_698;
  wire and_dcpl_700;
  wire or_tmp_238;
  wire or_tmp_242;
  wire and_dcpl_701;
  wire and_dcpl_707;
  wire or_dcpl_713;
  wire or_tmp_253;
  wire nor_tmp_135;
  wire nor_tmp_136;
  wire mux_tmp_211;
  wire mux_tmp_215;
  wire or_tmp_265;
  wire and_dcpl_711;
  wire and_dcpl_713;
  wire or_tmp_268;
  wire or_tmp_270;
  wire mux_tmp_220;
  wire or_tmp_275;
  wire mux_tmp_225;
  wire and_dcpl_714;
  wire mux_tmp_233;
  wire mux_tmp_237;
  wire or_tmp_294;
  wire mux_tmp_238;
  wire and_dcpl_721;
  wire or_tmp_298;
  wire mux_tmp_241;
  wire nor_tmp_159;
  wire or_tmp_300;
  wire mux_tmp_242;
  wire mux_tmp_247;
  wire mux_tmp_250;
  wire or_tmp_307;
  wire mux_tmp_259;
  wire or_tmp_315;
  wire mux_tmp_260;
  wire or_tmp_317;
  wire mux_tmp_262;
  wire mux_tmp_264;
  wire mux_tmp_266;
  wire or_tmp_329;
  wire or_tmp_338;
  wire mux_tmp_279;
  wire or_tmp_345;
  wire and_dcpl_725;
  wire and_dcpl_726;
  wire or_dcpl_715;
  wire and_dcpl_727;
  wire nor_tmp_197;
  wire nor_tmp_199;
  wire and_dcpl_728;
  wire and_dcpl_731;
  wire not_tmp_456;
  wire or_tmp_353;
  wire not_tmp_457;
  wire and_dcpl_732;
  wire and_dcpl_738;
  wire or_tmp_360;
  wire mux_tmp_295;
  wire mux_tmp_296;
  wire mux_tmp_301;
  wire mux_tmp_304;
  wire or_tmp_369;
  wire or_tmp_377;
  wire mux_tmp_312;
  wire or_tmp_391;
  wire mux_tmp_320;
  wire or_tmp_399;
  wire mux_tmp_327;
  wire or_tmp_406;
  wire and_dcpl_742;
  wire or_tmp_418;
  wire or_dcpl_717;
  wire [3:0] pe_config_manager_counter_sva_mx1;
  wire [4:0] operator_4_false_acc_sdt_sva_1;
  wire [5:0] nl_operator_4_false_acc_sdt_sva_1;
  reg [3:0] pe_config_num_manager_sva;
  wire state_0_sva_mx1;
  wire while_if_and_tmp_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiWrite_switch_lp_nor_tmp_1;
  reg pe_config_is_valid_sva;
  reg pe_config_is_zero_first_sva;
  reg pe_manager_zero_active_sva;
  reg pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  reg pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  reg PECore_UpdateFSM_switch_lp_and_7_itm_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
  reg PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  reg [8:0] operator_8_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_8_false_acc_sdt_sva_1;
  wire PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  wire PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1;
  reg PECore_RunFSM_switch_lp_nor_tmp_1;
  reg [1:0] state_2_1_sva;
  reg state_0_sva;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0;
  reg PECore_RunFSM_switch_lp_equal_tmp_1_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  reg weight_mem_run_3_for_land_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg input_read_req_valid_lpi_1_dfm_1_11;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9;
  reg rva_in_reg_rw_sva_11;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_11;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_11;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_11;
  wire PECore_RunScale_if_for_1_operator_32_true_slc_32_1_svs_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_11;
  wire PECore_RunScale_if_for_2_operator_32_true_slc_32_1_svs_1;
  wire PECore_RunScale_if_for_3_operator_32_true_slc_32_1_svs_1;
  wire PECore_RunScale_if_for_4_operator_32_true_slc_32_1_svs_1;
  wire PECore_RunScale_if_for_5_operator_32_true_slc_32_1_svs_1;
  wire PECore_RunScale_if_for_6_operator_32_true_slc_32_1_svs_1;
  wire PECore_RunScale_if_for_7_operator_32_true_slc_32_1_svs_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_11;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  wire PECore_UpdateFSM_switch_lp_equal_tmp_6;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  wire PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
  wire PECore_UpdateFSM_switch_lp_nor_tmp_1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
  wire [7:0] pe_config_input_counter_sva_mx1;
  wire [8:0] operator_16_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_16_false_acc_sdt_sva_1;
  reg [7:0] pe_manager_num_input_sva;
  reg [7:0] pe_config_num_output_sva;
  wire PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8;
  reg weight_mem_run_3_for_land_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  wire PECore_RunScale_if_for_8_operator_32_true_slc_32_1_svs_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_10;
  wire PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  reg PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
  wire weight_mem_run_3_for_land_lpi_1_dfm_1_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_380_itm_1;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_363_itm_1;
  wire weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  wire weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_359_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_153_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_141_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_5_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_4_itm_1;
  wire weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_127_sva_1;
  reg input_write_req_valid_lpi_1_dfm_1_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1;
  wire input_write_req_valid_lpi_1_dfm_5;
  wire input_mem_banks_write_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1;
  reg [14:0] pe_manager_base_input_sva;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1;
  reg rva_in_reg_rw_sva_5;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_4;
  wire PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3;
  reg rva_in_reg_rw_sva_st_1_11;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11;
  reg while_stage_0_13;
  reg input_read_req_valid_lpi_1_dfm_1_10;
  reg rva_in_reg_rw_sva_10;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8;
  reg rva_in_reg_rw_sva_st_1_10;
  reg rva_in_reg_rw_sva_st_10;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_10;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_10;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_9;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9;
  reg while_stage_0_11;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  reg while_stage_0_10;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  reg while_stage_0_9;
  reg rva_in_reg_rw_sva_st_1_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  reg rva_in_reg_rw_sva_st_1_5;
  reg while_stage_0_7;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_1;
  reg while_stage_0_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1;
  reg while_stage_0_5;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0;
  reg while_stage_0_4;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  reg while_stage_0_3;
  reg PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  reg [1:0] state_2_1_sva_dfm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_9;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
  reg while_stage_0_8;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_1;
  reg rva_in_reg_rw_sva_st_1_4;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_2;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  reg rva_in_reg_rw_sva_st_9;
  reg input_read_req_valid_lpi_1_dfm_1_9;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
  reg rva_in_reg_rw_sva_st_1_9;
  reg rva_in_reg_rw_sva_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1;
  reg rva_in_reg_rw_sva_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1;
  reg rva_in_reg_rw_sva_st_8;
  reg input_read_req_valid_lpi_1_dfm_1_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  reg rva_in_reg_rw_sva_st_1_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  reg rva_in_reg_rw_sva_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
  reg rva_in_reg_rw_sva_st_7;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  reg input_read_req_valid_lpi_1_dfm_1_7;
  reg rva_in_reg_rw_sva_st_1_7;
  reg rva_in_reg_rw_sva_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
  reg rva_in_reg_rw_sva_st_6;
  reg input_read_req_valid_lpi_1_dfm_1_6;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
  reg rva_in_reg_rw_sva_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
  reg rva_in_reg_rw_sva_st_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
  reg rva_in_reg_rw_sva_3;
  reg rva_in_reg_rw_sva_st_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2;
  reg input_read_req_valid_lpi_1_dfm_1_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
  reg input_read_req_valid_lpi_1_dfm_1_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
  reg input_read_req_valid_lpi_1_dfm_1_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1;
  reg [3:0] while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_10;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_10;
  reg while_stage_0_12;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_336_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_328_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_11;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_2;
  reg while_and_1282_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_4_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_1_sva;
  reg [7:0] weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_3_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_2_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_1_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_6_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_0_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_3_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs;
  wire operator_7_false_1_operator_7_false_1_or_mdf_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_1_sva_1;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_3_2_0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_3_2_0;
  reg [14:0] weight_read_addrs_7_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_5_lpi_1_dfm_1;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_2_2_0;
  reg [14:0] pe_manager_base_weight_sva;
  reg [14:0] weight_read_addrs_3_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_1_lpi_1_dfm_1;
  wire [3:0] pe_manager_base_weight_sva_mx1_3_0;
  wire pe_manager_base_weight_sva_mx3_0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  wire [11:0] nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1;
  reg [7:0] while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4;
  wire [7:0] input_write_addrs_lpi_1_dfm_2;
  wire [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_2;
  wire PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
  wire while_and_234_rgt;
  wire while_and_238_rgt;
  wire while_and_242_rgt;
  wire while_and_246_rgt;
  wire while_and_250_rgt;
  wire while_and_254_rgt;
  wire while_and_258_rgt;
  wire while_and_262_rgt;
  wire while_and_266_rgt;
  wire while_and_270_rgt;
  wire while_and_274_rgt;
  wire while_and_278_rgt;
  wire while_and_282_rgt;
  wire while_and_286_rgt;
  wire while_and_290_rgt;
  wire while_and_294_rgt;
  wire while_and_298_rgt;
  wire while_and_302_rgt;
  wire while_and_306_rgt;
  wire while_and_310_rgt;
  wire while_and_314_rgt;
  wire while_and_318_rgt;
  wire while_and_322_rgt;
  wire while_and_326_rgt;
  wire while_and_330_rgt;
  wire while_and_334_rgt;
  wire while_and_338_rgt;
  wire while_and_342_rgt;
  wire while_and_346_rgt;
  wire while_and_350_rgt;
  wire while_and_354_rgt;
  wire while_and_358_rgt;
  wire while_and_362_rgt;
  wire while_and_366_rgt;
  wire while_and_370_rgt;
  wire while_and_374_rgt;
  wire while_and_378_rgt;
  wire while_and_382_rgt;
  wire while_and_386_rgt;
  wire while_and_390_rgt;
  wire while_and_394_rgt;
  wire while_and_398_rgt;
  wire while_and_402_rgt;
  wire while_and_406_rgt;
  wire while_and_410_rgt;
  wire while_and_414_rgt;
  wire while_and_418_rgt;
  wire while_and_422_rgt;
  wire while_and_426_rgt;
  wire while_and_430_rgt;
  wire while_and_434_rgt;
  wire while_and_438_rgt;
  wire while_and_442_rgt;
  wire while_and_446_rgt;
  wire while_and_450_rgt;
  wire while_and_454_rgt;
  wire while_and_458_rgt;
  wire while_and_462_rgt;
  wire while_and_466_rgt;
  wire while_and_470_rgt;
  wire while_and_474_rgt;
  wire while_and_478_rgt;
  wire while_and_482_rgt;
  wire while_and_486_rgt;
  wire while_and_490_rgt;
  wire while_and_494_rgt;
  wire while_and_498_rgt;
  wire while_and_502_rgt;
  wire while_and_506_rgt;
  wire while_and_510_rgt;
  wire while_and_514_rgt;
  wire while_and_518_rgt;
  wire while_and_522_rgt;
  wire while_and_526_rgt;
  wire while_and_530_rgt;
  wire while_and_534_rgt;
  wire while_and_538_rgt;
  wire while_and_542_rgt;
  wire while_and_546_rgt;
  wire while_and_550_rgt;
  wire while_and_554_rgt;
  wire while_and_558_rgt;
  wire while_and_562_rgt;
  wire while_and_566_rgt;
  wire while_and_570_rgt;
  wire while_and_574_rgt;
  wire while_and_578_rgt;
  wire while_and_582_rgt;
  wire while_and_586_rgt;
  wire while_and_590_rgt;
  wire while_and_594_rgt;
  wire while_and_598_rgt;
  wire while_and_602_rgt;
  wire while_and_606_rgt;
  wire while_and_610_rgt;
  wire while_and_614_rgt;
  wire while_and_618_rgt;
  wire while_and_622_rgt;
  wire while_and_626_rgt;
  wire while_and_630_rgt;
  wire while_and_634_rgt;
  wire while_and_638_rgt;
  wire while_and_642_rgt;
  wire while_and_646_rgt;
  wire while_and_650_rgt;
  wire while_and_654_rgt;
  wire while_and_658_rgt;
  wire while_and_662_rgt;
  wire while_and_666_rgt;
  wire while_and_670_rgt;
  wire while_and_674_rgt;
  wire while_and_678_rgt;
  wire while_and_682_rgt;
  wire while_and_686_rgt;
  wire while_and_690_rgt;
  wire while_and_694_rgt;
  wire while_and_698_rgt;
  wire while_and_702_rgt;
  wire while_and_706_rgt;
  wire while_and_710_rgt;
  wire while_and_714_rgt;
  wire while_and_718_rgt;
  wire while_and_722_rgt;
  wire while_and_726_rgt;
  wire while_and_730_rgt;
  wire while_and_734_rgt;
  wire while_and_738_rgt;
  wire while_and_742_rgt;
  wire while_and_746_rgt;
  wire while_and_750_rgt;
  wire while_and_754_rgt;
  wire while_and_758_rgt;
  wire while_and_762_rgt;
  wire while_and_766_rgt;
  wire while_and_770_rgt;
  wire while_and_774_rgt;
  wire while_and_778_rgt;
  wire while_and_782_rgt;
  wire while_and_786_rgt;
  wire while_and_790_rgt;
  wire while_and_794_rgt;
  wire while_and_798_rgt;
  wire while_and_802_rgt;
  wire while_and_806_rgt;
  wire while_and_810_rgt;
  wire while_and_814_rgt;
  wire while_and_818_rgt;
  wire while_and_822_rgt;
  wire while_and_826_rgt;
  wire while_and_830_rgt;
  wire while_and_834_rgt;
  wire while_and_838_rgt;
  wire while_and_842_rgt;
  wire while_and_846_rgt;
  wire while_and_850_rgt;
  wire while_and_854_rgt;
  wire while_and_858_rgt;
  wire while_and_862_rgt;
  wire while_and_866_rgt;
  wire while_and_870_rgt;
  wire while_and_874_rgt;
  wire while_and_878_rgt;
  wire while_and_882_rgt;
  wire while_and_886_rgt;
  wire while_and_890_rgt;
  wire while_and_894_rgt;
  wire while_and_898_rgt;
  wire while_and_902_rgt;
  wire while_and_906_rgt;
  wire while_and_910_rgt;
  wire while_and_914_rgt;
  wire while_and_918_rgt;
  wire while_and_922_rgt;
  wire while_and_926_rgt;
  wire while_and_930_rgt;
  wire while_and_934_rgt;
  wire while_and_938_rgt;
  wire while_and_942_rgt;
  wire while_and_946_rgt;
  wire while_and_950_rgt;
  wire while_and_954_rgt;
  wire while_and_958_rgt;
  wire while_and_962_rgt;
  wire while_and_966_rgt;
  wire while_and_970_rgt;
  wire while_and_974_rgt;
  wire while_and_978_rgt;
  wire while_and_982_rgt;
  wire while_and_986_rgt;
  wire while_and_990_rgt;
  wire while_and_994_rgt;
  wire while_and_998_rgt;
  wire while_and_1002_rgt;
  wire while_and_1006_rgt;
  wire while_and_1010_rgt;
  wire while_and_1014_rgt;
  wire while_and_1018_rgt;
  wire while_and_1022_rgt;
  wire while_and_1026_rgt;
  wire while_and_1030_rgt;
  wire while_and_1034_rgt;
  wire while_and_1038_rgt;
  wire while_and_1042_rgt;
  wire while_and_1046_rgt;
  wire while_and_1050_rgt;
  wire while_and_1054_rgt;
  wire while_and_1058_rgt;
  wire while_and_1062_rgt;
  wire while_and_1066_rgt;
  wire while_and_1070_rgt;
  wire while_and_1074_rgt;
  wire while_and_1078_rgt;
  wire while_and_1082_rgt;
  wire while_and_1086_rgt;
  wire while_and_1090_rgt;
  wire while_and_1094_rgt;
  wire while_and_1098_rgt;
  wire while_and_1102_rgt;
  wire while_and_1106_rgt;
  wire while_and_1110_rgt;
  wire while_and_1114_rgt;
  wire while_and_1118_rgt;
  wire while_and_1122_rgt;
  wire while_and_1126_rgt;
  wire while_and_1130_rgt;
  wire while_and_1134_rgt;
  wire while_and_1138_rgt;
  wire while_and_1142_rgt;
  wire while_and_1146_rgt;
  wire while_and_1150_rgt;
  wire while_and_1154_rgt;
  wire while_and_1158_rgt;
  wire while_and_1162_rgt;
  wire while_and_1166_rgt;
  wire while_and_1170_rgt;
  wire while_and_1174_rgt;
  wire while_and_1178_rgt;
  wire while_and_1182_rgt;
  wire while_and_1186_rgt;
  wire while_and_1190_rgt;
  wire while_and_1194_rgt;
  wire while_and_1198_rgt;
  wire while_and_1202_rgt;
  wire while_and_1206_rgt;
  wire while_and_1210_rgt;
  wire while_and_1214_rgt;
  wire while_and_1218_rgt;
  wire while_and_1222_rgt;
  wire while_and_1226_rgt;
  wire while_and_1230_rgt;
  wire while_and_1234_rgt;
  wire while_and_1238_rgt;
  wire while_and_1242_rgt;
  wire while_and_1246_rgt;
  wire while_and_1250_rgt;
  wire while_and_1254_rgt;
  wire weight_mem_banks_read_1_for_mux_cse;
  wire weight_mem_banks_read_1_for_mux_1_cse;
  wire weight_mem_banks_read_1_for_mux_4_cse;
  wire weight_mem_banks_read_1_for_mux_5_cse;
  wire weight_mem_banks_read_1_for_mux_8_cse;
  wire weight_mem_banks_read_1_for_mux_9_cse;
  wire weight_mem_banks_read_1_for_mux_12_cse;
  wire weight_mem_banks_read_1_for_mux_13_cse;
  wire weight_mem_banks_read_1_for_mux_16_cse;
  wire weight_mem_banks_read_1_for_mux_17_cse;
  wire weight_mem_banks_read_1_for_mux_20_cse;
  wire weight_mem_banks_read_1_for_mux_21_cse;
  wire weight_mem_banks_read_1_for_mux_24_cse;
  wire weight_mem_banks_read_1_for_mux_25_cse;
  wire weight_mem_banks_read_1_for_mux_28_cse;
  wire weight_mem_banks_read_1_for_mux_29_cse;
  wire weight_mem_banks_write_if_for_if_mux_8_cse;
  wire weight_mem_banks_write_if_for_if_mux_9_cse;
  wire weight_mem_banks_read_for_mux_cse;
  wire weight_mem_banks_read_for_mux_1_cse;
  wire weight_mem_banks_write_if_for_if_mux_12_cse;
  wire weight_mem_banks_write_if_for_if_mux_13_cse;
  wire weight_mem_banks_read_for_mux_4_cse;
  wire weight_mem_banks_read_for_mux_5_cse;
  wire weight_mem_banks_write_if_for_if_mux_16_cse;
  wire weight_mem_banks_write_if_for_if_mux_17_cse;
  wire weight_mem_banks_read_for_mux_8_cse;
  wire weight_mem_banks_read_for_mux_9_cse;
  wire weight_mem_banks_write_if_for_if_mux_20_cse;
  wire weight_mem_banks_write_if_for_if_mux_21_cse;
  wire weight_mem_banks_read_for_mux_12_cse;
  wire weight_mem_banks_read_for_mux_13_cse;
  wire weight_mem_banks_write_if_for_if_mux_24_cse;
  wire weight_mem_banks_write_if_for_if_mux_25_cse;
  wire weight_mem_banks_read_for_mux_16_cse;
  wire weight_mem_banks_read_for_mux_17_cse;
  wire weight_mem_banks_write_if_for_if_mux_28_cse;
  wire weight_mem_banks_write_if_for_if_mux_29_cse;
  wire weight_mem_banks_read_for_mux_20_cse;
  wire weight_mem_banks_read_for_mux_21_cse;
  wire weight_mem_banks_write_if_for_if_mux_32_cse;
  wire weight_mem_banks_write_if_for_if_mux_33_cse;
  wire weight_mem_banks_read_for_mux_24_cse;
  wire weight_mem_banks_read_for_mux_25_cse;
  wire weight_mem_banks_write_if_for_if_mux_36_cse;
  wire weight_mem_banks_write_if_for_if_mux_37_cse;
  wire weight_mem_banks_read_for_mux_28_cse;
  wire weight_mem_banks_read_for_mux_29_cse;
  wire input_mem_banks_write_1_if_for_if_mux_cse;
  wire input_mem_banks_write_1_if_for_if_mux_1_cse;
  wire input_mem_banks_read_1_for_mux_cse;
  wire input_mem_banks_read_1_for_mux_1_cse;
  wire input_mem_banks_write_if_for_if_mux_cse;
  wire input_mem_banks_write_if_for_if_mux_1_cse;
  wire input_mem_banks_read_for_mux_cse;
  wire input_mem_banks_read_for_mux_1_cse;
  reg reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_63_cse;
  reg reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_40_cse;
  reg reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_7_cse;
  reg reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_1_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_act_port_Push_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire rva_out_reg_data_and_cse;
  wire accum_vector_data_and_cse;
  wire weight_port_read_out_data_and_1_cse;
  wire weight_port_read_out_data_and_16_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_cse;
  reg reg_rva_in_reg_rw_sva_st_1_1_cse;
  wire or_142_cse;
  wire weight_port_read_out_data_and_50_cse;
  wire weight_port_read_out_data_and_78_cse;
  wire weight_port_read_out_data_and_109_cse;
  reg reg_weight_mem_run_3_for_5_and_15_itm_1_cse;
  reg reg_weight_mem_run_3_for_5_and_16_itm_1_cse;
  reg reg_weight_mem_run_3_for_5_and_6_itm_1_cse;
  wire or_188_cse;
  wire operator_15_false_1_and_cse;
  wire pe_config_num_manager_and_cse;
  wire PECore_DecodeAxiWrite_switch_lp_and_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
  reg [2:0] reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
  wire pe_manager_num_input_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_or_3_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_36_cse;
  wire Arbiter_8U_Roundrobin_pick_and_26_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_24_cse;
  wire Arbiter_8U_Roundrobin_pick_and_20_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_10_cse;
  wire Arbiter_8U_Roundrobin_pick_and_13_cse;
  wire or_185_cse;
  wire [1:0] state_mux_1_cse;
  wire and_279_cse;
  wire and_572_cse;
  wire and_576_cse;
  wire and_542_cse;
  wire and_537_cse;
  wire and_626_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_7_or_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  wire while_and_21_cse;
  wire or_50_cse;
  wire while_and_45_cse;
  wire nor_279_cse;
  wire nor_276_cse;
  wire nor_280_cse;
  wire nor_284_cse;
  wire nand_35_cse;
  wire nor_335_cse;
  wire while_and_1256_cse;
  wire while_while_nor_259_cse;
  wire and_777_cse;
  wire and_779_cse;
  wire and_782_cse;
  wire and_784_cse;
  wire and_783_cse;
  wire and_778_cse;
  wire and_788_cse;
  wire and_790_cse;
  wire and_789_cse;
  wire and_780_cse;
  wire and_810_cse;
  wire and_814_cse;
  wire and_815_cse;
  wire and_825_cse;
  wire and_818_cse;
  wire and_819_cse;
  wire and_816_cse;
  wire and_820_cse;
  wire and_843_cse;
  wire and_844_cse;
  wire and_997_cse;
  wire and_999_cse;
  wire and_996_cse;
  wire and_858_cse;
  wire and_998_cse;
  wire and_857_cse;
  wire and_869_cse;
  wire and_867_cse;
  wire and_873_cse;
  wire and_875_cse;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_82_cse;
  wire nor_423_cse;
  wire nand_62_cse;
  wire and_893_cse;
  wire and_900_cse;
  wire and_898_cse;
  wire and_897_cse;
  wire and_899_cse;
  wire and_890_cse;
  wire and_905_cse;
  wire and_907_cse;
  wire and_910_cse;
  wire and_915_cse;
  wire and_906_cse;
  wire and_1000_cse;
  wire and_1001_cse;
  wire and_1007_cse;
  wire and_1008_cse;
  wire and_1009_cse;
  wire and_1002_cse;
  wire and_1004_cse;
  wire and_1003_cse;
  wire and_1006_cse;
  wire and_937_cse;
  wire and_944_cse;
  wire and_943_cse;
  wire and_945_cse;
  wire and_936_cse;
  wire and_1005_cse;
  wire and_958_cse;
  reg Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2;
  wire while_if_and_2_m1c;
  wire weight_mem_run_3_for_5_and_163_cse;
  wire weight_mem_run_3_for_5_and_162_cse;
  wire mux_115_cse;
  wire pe_config_is_valid_and_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_12_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_55_cse;
  wire Arbiter_8U_Roundrobin_pick_and_44_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_63_cse;
  wire Arbiter_8U_Roundrobin_pick_and_52_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_85_cse;
  wire Arbiter_8U_Roundrobin_pick_and_74_cse;
  wire and_352_cse;
  wire pe_config_input_counter_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse;
  wire and_115_cse;
  wire and_122_cse;
  wire or_944_cse;
  wire or_945_cse;
  wire or_1079_cse;
  wire or_1140_cse;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1;
  wire PECore_DecodeAxiWrite_switch_lp_or_5_cse_1;
  wire Arbiter_8U_Roundrobin_pick_and_14_cse;
  wire Arbiter_8U_Roundrobin_pick_and_8_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse;
  wire mux_192_cse;
  wire mux_335_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0;
  wire and_570_rmff;
  wire and_567_rmff;
  wire and_564_rmff;
  wire and_561_rmff;
  wire and_558_rmff;
  wire and_555_rmff;
  wire and_551_rmff;
  wire and_548_rmff;
  wire and_541_rmff;
  wire and_544_rmff;
  wire and_535_rmff;
  wire and_538_rmff;
  wire and_574_rmff;
  reg [35:0] accum_vector_data_0_35_0_sva;
  reg [35:0] accum_vector_data_7_35_0_sva;
  reg [35:0] accum_vector_data_6_35_0_sva;
  reg [35:0] accum_vector_data_5_35_0_sva;
  reg [35:0] accum_vector_data_4_35_0_sva;
  reg [35:0] accum_vector_data_3_35_0_sva;
  reg [35:0] accum_vector_data_2_35_0_sva;
  reg [35:0] accum_vector_data_1_35_0_sva;
  reg [7:0] pe_config_output_counter_sva;
  reg [7:0] pe_config_input_counter_sva;
  reg [31:0] act_port_reg_data_255_224_sva_dfm_1_1;
  wire [31:0] act_port_reg_data_223_192_sva_dfm_3;
  wire [31:0] act_port_reg_data_191_160_sva_dfm_3;
  wire [31:0] act_port_reg_data_159_128_sva_dfm_3;
  wire [31:0] act_port_reg_data_127_96_sva_dfm_3;
  wire [31:0] act_port_reg_data_95_64_sva_dfm_3;
  wire [31:0] act_port_reg_data_63_32_sva_dfm_3;
  wire [31:0] act_port_reg_data_31_0_sva_dfm_3;
  reg [15:0] rva_out_reg_data_255_240_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_239_224_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_223_208_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_207_192_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_191_176_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_175_160_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_159_144_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_143_128_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_6;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_6;
  reg rva_out_reg_data_63_sva_dfm_4_6;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_6;
  reg rva_out_reg_data_47_sva_dfm_4_6;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_6;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_6;
  wire rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_31_mx0;
  wire rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_24_mx0;
  wire [6:0] rva_out_reg_data_23_17_sva_dfm_7;
  wire rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_16_mx0;
  wire [6:0] rva_out_reg_data_15_9_sva_dfm_7;
  wire rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_8_mx0;
  wire [6:0] rva_out_reg_data_7_1_sva_dfm_7;
  wire rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_0_mx0;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_4;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0;
  reg weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
  reg [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1;
  reg [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1;
  reg [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1;
  reg weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  reg [15:0] weight_port_read_out_data_3_15_sva_dfm_1;
  reg [255:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_5;
  reg [15:0] weight_mem_run_3_for_5_mux_62_itm_1;
  reg [255:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
  reg [15:0] weight_port_read_out_data_0_0_sva_dfm_1_1;
  reg [15:0] weight_port_read_out_data_0_3_sva_dfm_1_1;
  reg [15:0] weight_port_read_out_data_0_2_sva_dfm_1_1;
  reg [15:0] weight_mem_run_3_for_5_mux_5_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_4_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_7_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_6_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_9_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_8_itm_1;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_1;
  reg [15:0] weight_mem_run_3_for_5_mux_13_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_12_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_15_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_14_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_97_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_96_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_99_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_98_itm_1;
  reg [15:0] rva_out_reg_data_143_128_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_175_160_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_159_144_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_207_192_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_191_176_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_239_224_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_223_208_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_1;
  reg [15:0] rva_out_reg_data_255_240_sva_dfm_4_1;
  reg [15:0] weight_mem_run_3_for_5_mux_111_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_110_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_17_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_16_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_19_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_18_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_21_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_20_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_23_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_22_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_25_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_24_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_27_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_26_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_29_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_28_itm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  reg [15:0] weight_port_read_out_data_1_15_sva_dfm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_30_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_81_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_80_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_83_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_82_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_85_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_84_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_87_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_86_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_89_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_88_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_91_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_90_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_93_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_92_itm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  reg [15:0] weight_port_read_out_data_2_1_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
  reg [15:0] weight_port_read_out_data_2_0_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
  reg [15:0] weight_port_read_out_data_2_3_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
  reg [15:0] weight_port_read_out_data_2_2_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
  reg [15:0] weight_port_read_out_data_2_5_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
  reg [15:0] weight_port_read_out_data_2_4_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
  reg [15:0] weight_port_read_out_data_2_7_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
  reg [15:0] weight_port_read_out_data_2_6_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
  reg [15:0] weight_port_read_out_data_2_9_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
  reg [15:0] weight_port_read_out_data_2_8_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
  reg [15:0] weight_port_read_out_data_2_11_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
  reg [15:0] weight_port_read_out_data_2_10_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
  reg [15:0] weight_port_read_out_data_2_13_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
  reg [15:0] weight_port_read_out_data_2_12_sva_dfm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_47_itm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014;
  reg [15:0] weight_port_read_out_data_2_14_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  reg [15:0] weight_port_read_out_data_4_1_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
  reg [15:0] weight_port_read_out_data_4_0_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
  reg [15:0] weight_port_read_out_data_4_3_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
  reg [15:0] weight_port_read_out_data_4_2_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
  reg [15:0] weight_port_read_out_data_4_5_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
  reg [15:0] weight_port_read_out_data_4_4_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
  reg [15:0] weight_port_read_out_data_4_7_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
  reg [15:0] weight_port_read_out_data_4_6_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
  reg [15:0] weight_port_read_out_data_4_9_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
  reg [15:0] weight_port_read_out_data_4_8_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
  reg [15:0] weight_port_read_out_data_4_11_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
  reg [15:0] weight_port_read_out_data_4_10_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
  reg [15:0] weight_port_read_out_data_4_13_sva_dfm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
  reg [15:0] weight_port_read_out_data_4_12_sva_dfm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_79_itm_1;
  reg [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014;
  reg [15:0] weight_port_read_out_data_4_14_sva_dfm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_49_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_48_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_51_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_50_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_53_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_52_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_55_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_54_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_57_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_56_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_59_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_58_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_61_itm_1;
  reg [15:0] weight_mem_run_3_for_5_mux_60_itm_1;
  reg [15:0] weight_write_data_data_0_15_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_14_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_13_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_12_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_11_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_10_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_9_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_8_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
  reg [15:0] weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
  reg [14:0] weight_write_addrs_lpi_1_dfm_1_2;
  reg [15:0] weight_write_data_data_0_15_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_14_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_13_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_12_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_11_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_10_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_9_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_8_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_7_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_6_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_5_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_4_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_3_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_2_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_1_lpi_1_dfm_1_3_2;
  reg [15:0] weight_write_data_data_0_0_lpi_1_dfm_1_3_2;
  reg [11:0] weight_write_addrs_lpi_1_dfm_1_3_14_3;
  wire and_dcpl_743;
  wire or_dcpl;
  wire or_dcpl_719;
  wire or_dcpl_720;
  reg [255:0] input_mem_banks_read_read_data_lpi_1_dfm_1_4;
  reg [255:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1;
  reg [255:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1;
  reg [255:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1;
  reg [255:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1;
  wire [255:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0;
  wire [239:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0;
  reg [1:0] weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_itm_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_231_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_28;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1;
  wire and_1025_cse;
  wire and_1026_cse;
  wire and_1027_cse;
  wire and_1017_cse;
  wire and_1018_cse;
  wire and_1019_cse;
  wire and_1020_cse;
  wire and_1021_cse;
  wire and_1022_cse;
  wire nor_472_cse;
  wire and_1038_cse;
  wire and_1039_cse;
  wire and_1040_cse;
  wire and_1041_cse;
  wire and_1042_cse;
  wire nor_473_cse;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1;
  wire [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm;
  wire mux_129_itm;
  wire mux_136_itm;
  wire mux_158_itm;
  wire mux_172_itm;
  wire mux_257_itm;
  wire mux_276_itm;
  wire mux_311_itm;
  wire mux_324_itm;
  reg weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  reg [15:0] weight_port_read_out_data_0_3_sva;
  reg [15:0] weight_port_read_out_data_0_2_sva;
  reg [14:0] pe_manager_base_bias_sva;
  reg pe_config_is_cluster_sva;
  reg pe_config_is_bias_sva;
  reg [3:0] pe_config_manager_counter_sva;
  reg [31:0] act_port_reg_data_127_96_sva;
  reg [31:0] act_port_reg_data_159_128_sva;
  reg [31:0] act_port_reg_data_95_64_sva;
  reg [31:0] act_port_reg_data_191_160_sva;
  reg [31:0] act_port_reg_data_63_32_sva;
  reg [31:0] act_port_reg_data_223_192_sva;
  reg [31:0] act_port_reg_data_31_0_sva;
  reg [31:0] act_port_reg_data_255_224_sva;
  reg [15:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8;
  reg [255:0] input_mem_banks_bank_a_0_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_1_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_2_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_3_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_4_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_5_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_6_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_7_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_8_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_9_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_10_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_11_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_12_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_13_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_14_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_15_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_16_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_17_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_18_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_19_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_20_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_21_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_22_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_23_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_24_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_25_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_26_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_27_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_28_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_29_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_30_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_31_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_32_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_33_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_34_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_35_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_36_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_37_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_38_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_39_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_40_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_41_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_42_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_43_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_44_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_45_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_46_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_47_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_48_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_49_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_50_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_51_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_52_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_53_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_54_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_55_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_56_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_57_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_58_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_59_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_60_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_61_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_62_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_63_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_64_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_65_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_66_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_67_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_68_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_69_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_70_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_71_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_72_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_73_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_74_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_75_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_76_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_77_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_78_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_79_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_80_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_81_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_82_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_83_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_84_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_85_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_86_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_87_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_88_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_89_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_90_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_91_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_92_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_93_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_94_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_95_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_96_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_97_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_98_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_99_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_100_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_101_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_102_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_103_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_104_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_105_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_106_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_107_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_108_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_109_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_110_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_111_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_112_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_113_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_114_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_115_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_116_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_117_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_118_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_119_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_120_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_121_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_122_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_123_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_124_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_125_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_126_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_127_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_128_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_129_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_130_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_131_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_132_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_133_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_134_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_135_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_136_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_137_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_138_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_139_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_140_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_141_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_142_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_143_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_144_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_145_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_146_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_147_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_148_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_149_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_150_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_151_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_152_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_153_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_154_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_155_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_156_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_157_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_158_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_159_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_160_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_161_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_162_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_163_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_164_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_165_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_166_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_167_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_168_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_169_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_170_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_171_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_172_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_173_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_174_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_175_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_176_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_177_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_178_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_179_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_180_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_181_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_182_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_183_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_184_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_185_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_186_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_187_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_188_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_189_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_190_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_191_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_192_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_193_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_194_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_195_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_196_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_197_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_198_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_199_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_200_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_201_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_202_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_203_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_204_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_205_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_206_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_207_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_208_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_209_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_210_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_211_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_212_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_213_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_214_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_215_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_216_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_217_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_218_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_219_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_220_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_221_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_222_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_223_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_224_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_225_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_226_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_227_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_228_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_229_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_230_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_231_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_232_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_233_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_234_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_235_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_236_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_237_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_238_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_239_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_240_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_241_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_242_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_243_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_244_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_245_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_246_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_247_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_248_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_249_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_250_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_251_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_252_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_253_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_254_sva_dfm_2;
  reg [255:0] input_mem_banks_bank_a_255_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_0_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_4_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_5_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_6_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_7_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_8_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_9_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_10_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_11_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_12_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_13_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_14_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_0_15_sva_dfm_2;
  reg [15:0] weight_port_read_out_data_1_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_8_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_9_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_10_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_11_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_12_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_13_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_1_14_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_2_15_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_8_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_9_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_10_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_11_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_12_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_13_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_3_14_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_4_15_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_8_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_9_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_10_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_11_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_12_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_13_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_14_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_5_15_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_8_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_9_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_10_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_11_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_12_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_13_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_14_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_6_15_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_0_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_1_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_4_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_5_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_6_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_7_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_8_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_9_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_10_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_11_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_12_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_13_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_14_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_7_15_sva_dfm_1;
  reg rva_out_reg_data_24_sva_dfm_6;
  reg rva_out_reg_data_31_sva_dfm_6;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_6;
  reg rva_out_reg_data_16_sva_dfm_6;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_6;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_6;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_6;
  reg rva_out_reg_data_8_sva_dfm_6;
  reg [6:0] rva_out_reg_data_7_1_sva_dfm_6;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_6;
  reg rva_out_reg_data_0_sva_dfm_6;
  reg [255:0] weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1;
  reg [255:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1;
  reg [255:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1;
  reg [255:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1;
  reg [255:0] weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1;
  reg [255:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1;
  reg [255:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1;
  reg [15:0] rva_out_reg_data_255_240_sva_dfm_6;
  reg [15:0] rva_out_reg_data_239_224_sva_dfm_6;
  reg [15:0] rva_out_reg_data_223_208_sva_dfm_6;
  reg [15:0] rva_out_reg_data_207_192_sva_dfm_6;
  reg [15:0] rva_out_reg_data_191_176_sva_dfm_6;
  reg [15:0] rva_out_reg_data_175_160_sva_dfm_6;
  reg [15:0] rva_out_reg_data_159_144_sva_dfm_6;
  reg [15:0] rva_out_reg_data_143_128_sva_dfm_6;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_6;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_6;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_6;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_6;
  reg rva_out_reg_data_63_sva_dfm_6;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2;
  reg [35:0] accum_vector_data_7_35_0_sva_dfm_1_1;
  reg [35:0] accum_vector_data_6_35_0_sva_dfm_1_1;
  reg [35:0] accum_vector_data_5_35_0_sva_dfm_1_1;
  reg [35:0] accum_vector_data_4_35_0_sva_dfm_1_1;
  reg [35:0] accum_vector_data_3_35_0_sva_dfm_1_1;
  reg [35:0] accum_vector_data_2_35_0_sva_dfm_1_1;
  reg [35:0] accum_vector_data_1_35_0_sva_dfm_1_1;
  reg [35:0] accum_vector_data_0_35_0_sva_dfm_1_1;
  reg [3:0] pe_config_manager_counter_sva_dfm_3_1;
  reg [7:0] input_read_addrs_sva_1_1;
  wire [8:0] nl_input_read_addrs_sva_1_1;
  reg rva_out_reg_data_63_sva_dfm_4_4;
  reg rva_out_reg_data_63_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_79_64_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_95_80_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_111_96_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_127_112_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_143_128_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_143_128_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_143_128_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_143_128_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_159_144_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_159_144_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_159_144_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_159_144_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_175_160_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_175_160_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_175_160_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_175_160_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_191_176_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_191_176_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_191_176_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_191_176_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_207_192_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_207_192_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_207_192_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_207_192_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_223_208_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_223_208_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_223_208_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_223_208_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_239_224_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_239_224_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_239_224_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_239_224_sva_dfm_4_5;
  reg [15:0] rva_out_reg_data_255_240_sva_dfm_4_2;
  reg [15:0] rva_out_reg_data_255_240_sva_dfm_4_3;
  reg [15:0] rva_out_reg_data_255_240_sva_dfm_4_4;
  reg [15:0] rva_out_reg_data_255_240_sva_dfm_4_5;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_1;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_2;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_3;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_4;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_4_5;
  reg rva_out_reg_data_47_sva_dfm_4_4;
  reg rva_out_reg_data_47_sva_dfm_4_5;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_3;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_4_5;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_1;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_2;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_4;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_4_5;
  reg [15:0] weight_port_read_out_data_0_3_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_0_2_sva_dfm_1;
  reg [15:0] weight_port_read_out_data_0_0_sva_dfm_2_1;
  reg [15:0] weight_port_read_out_data_0_0_sva_dfm_3;
  reg [15:0] weight_port_read_out_data_0_0_sva_dfm_4;
  reg [15:0] weight_port_read_out_data_0_0_sva_dfm_5;
  reg [15:0] weight_port_read_out_data_0_0_sva_dfm_6;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_1_2;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_1_3;
  reg [14:0] rva_out_reg_data_62_48_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_5;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_5;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_1;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_2;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_4;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_5;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_6_1;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_7_1;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_8;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_9;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_10;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_11;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_1;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_2;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_3;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_4;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_5;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_6_1;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_7_1;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_8;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_9;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_1;
  reg [7:0] pe_config_output_counter_sva_dfm_1;
  reg [7:0] pe_config_input_counter_sva_dfm_1;
  reg [255:0] rva_in_reg_data_sva_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
  reg [14:0] weight_write_addrs_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_0_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_1_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_2_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_3_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_4_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_5_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_6_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_7_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_8_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_9_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_10_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_11_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_12_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_13_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_14_lpi_1_dfm_1_1;
  reg [15:0] weight_write_data_data_0_15_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_2;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_1;
  reg [255:0] input_mem_banks_read_read_data_lpi_1_dfm_1_2;
  reg [255:0] input_mem_banks_read_read_data_lpi_1_dfm_1_3;
  reg [10:0] PEManager_15U_GetWeightAddr_else_acc_3_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  reg [255:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
  reg [255:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
  reg [255:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
  reg [33:0] Datapath_for_6_ProductSum_for_acc_1_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_11;
  reg [14:0] pe_manager_base_weight_sva_dfm_3_1;
  reg [14:0] pe_manager_base_input_sva_dfm_3_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_11;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_11;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_39_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_71_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_37_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_69_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_36_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_68_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1;
  reg [15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_31_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_6;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_6;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_6;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_6;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_6;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_6;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_6;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_6;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_6;
  reg [15:0] weight_mem_banks_load_store_1_for_3_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1;
  reg [15:0] weight_mem_banks_load_store_1_for_5_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_104_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_14_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_36_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_2;
  reg weight_mem_run_3_for_5_and_146_itm_1;
  reg weight_mem_run_3_for_5_and_147_itm_1;
  reg weight_mem_run_3_for_5_and_148_itm_1;
  reg weight_mem_run_3_for_5_and_149_itm_1;
  reg weight_mem_run_3_for_5_and_150_itm_1;
  reg weight_mem_run_3_for_5_and_150_itm_2;
  reg weight_mem_run_3_for_5_and_151_itm_1;
  reg weight_mem_run_3_for_5_and_151_itm_2;
  reg weight_mem_run_3_for_5_and_152_itm_1;
  reg weight_mem_run_3_for_5_and_7_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
  reg weight_mem_run_3_for_5_and_12_itm_1;
  reg weight_mem_run_3_for_5_and_14_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1;
  reg weight_mem_run_3_for_5_and_126_itm_1;
  reg weight_mem_run_3_for_5_and_126_itm_2;
  reg weight_mem_run_3_for_5_and_132_itm_1;
  reg weight_mem_run_3_for_5_and_135_itm_1;
  reg weight_mem_run_3_for_5_and_135_itm_2;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2;
  reg weight_mem_run_3_for_5_and_140_itm_1;
  reg weight_mem_run_3_for_5_and_140_itm_2;
  reg weight_mem_run_3_for_5_and_142_itm_1;
  reg weight_mem_run_3_for_5_and_143_itm_1;
  reg weight_mem_run_3_for_5_and_144_itm_1;
  reg [14:0] PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1;
  reg while_if_mux_27_itm_1;
  reg PECore_PushAxiRsp_mux_10_itm_1;
  reg PECore_PushAxiRsp_mux_26_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  reg [239:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_1_255_16;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_3_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0;
  wire [31:0] act_port_reg_data_255_224_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_0_0_sva_dfm_1_mx0w0;
  wire [15:0] weight_port_read_out_data_0_0_sva_dfm_mx0w1;
  wire PECore_PushAxiRsp_if_else_mux_26_mx0w2;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_278_itm_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0;
  wire weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
  wire [14:0] pe_manager_base_weight_sva_mx2;
  wire [14:0] weight_read_addrs_1_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_3_lpi_1_dfm_1_1;
  wire [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_5_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_7_lpi_1_dfm_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  wire [7:0] pe_config_output_counter_sva_mx1;
  wire pe_config_is_zero_first_sva_mx1;
  wire pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  wire [15:0] weight_port_read_out_data_0_3_sva_mx0;
  wire [15:0] weight_port_read_out_data_0_2_sva_mx0;
  wire [15:0] weight_port_read_out_data_0_3_sva_dfm_2;
  wire [15:0] weight_port_read_out_data_0_2_sva_dfm_2;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_40_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_mx0w0;
  wire [14:0] pe_manager_base_input_sva_mx1;
  wire PECore_PushAxiRsp_if_else_mux_10_mx0w2;
  wire [15:0] rva_out_reg_data_255_240_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_239_224_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_223_208_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_207_192_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_191_176_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_175_160_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_159_144_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_143_128_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_127_112_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_111_96_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_95_80_sva_dfm_4_mx0w0;
  wire [15:0] rva_out_reg_data_79_64_sva_dfm_4_mx0w0;
  wire [14:0] rva_out_reg_data_62_48_sva_dfm_6_mx1;
  wire [6:0] rva_out_reg_data_46_40_sva_dfm_6_mx1;
  wire [3:0] rva_out_reg_data_39_36_sva_dfm_6_mx1;
  wire PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  wire [15:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1;
  wire weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_4;
  wire while_and_1285_cse_1;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_239_2000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_223_2000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_207_1000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_191_1000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_63_48_sva_1;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_175_1000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_79_64_sva_1;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_159_1000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_95_80_sva_1;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_143_1000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_111_9000000;
  wire [15:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_127_1000000;
  wire rva_out_reg_data_63_sva_dfm_7;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
  wire PECore_PushAxiRsp_if_asn_83;
  wire PECore_PushAxiRsp_if_asn_85;
  wire PECore_PushAxiRsp_if_asn_87;
  wire PECore_RunMac_asn_23;
  wire weight_mem_run_3_for_5_asn_445;
  wire weight_mem_run_3_for_5_asn_447;
  wire weight_mem_run_3_for_5_asn_449;
  wire weight_mem_run_3_for_5_asn_451;
  wire weight_mem_run_3_for_5_asn_453;
  wire weight_mem_run_3_for_5_asn_455;
  wire weight_mem_run_3_for_5_asn_457;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_411;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_419;
  wire PECore_PushAxiRsp_if_asn_91;
  wire PECore_PushAxiRsp_if_asn_93;
  wire PECore_PushAxiRsp_if_asn_95;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367;
  wire weight_mem_run_3_for_5_and_153;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126;
  wire weight_mem_run_3_for_5_and_157;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_128;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0;
  wire [15:0] weight_port_read_out_data_5_14_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_5_15_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_14_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_15_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_12_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_13_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_10_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_11_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_8_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_9_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_6_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_7_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_4_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_5_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_2_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_3_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_0_sva_dfm_3;
  wire [15:0] weight_port_read_out_data_7_1_sva_dfm_3;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse;
  reg reg_rva_in_reg_rw_sva_2_cse;
  reg reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_12_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_14_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_7_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_146_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_147_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_148_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_149_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_152_itm_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse;
  wire weight_mem_banks_load_store_for_else_and_80_ssc;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_15;
  reg [14:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_1_4_3_2;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_1_4_1_0;
  wire rva_out_reg_data_and_168_ssc;
  reg [3:0] rva_out_reg_data_30_25_sva_dfm_2_5_2;
  reg [1:0] rva_out_reg_data_30_25_sva_dfm_2_1_0;
  reg weight_port_read_out_data_0_1_sva_dfm_1_15;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_1_14_0;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_1_5_3_2;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_1_5_1_0;
  reg [3:0] rva_out_reg_data_30_25_sva_dfm_3_5_2;
  reg [1:0] rva_out_reg_data_30_25_sva_dfm_3_1_0;
  reg weight_port_read_out_data_0_1_sva_dfm_2_rsp_0;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_2_rsp_1;
  reg [3:0] rva_out_reg_data_30_25_sva_dfm_4_rsp_0;
  reg [1:0] rva_out_reg_data_30_25_sva_dfm_4_rsp_1;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd;
  reg [14:0] reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1;
  wire rva_out_reg_data_and_108_ssc;
  reg [3:0] reg_rva_out_reg_data_30_25_sva_dfm_5_ftd;
  reg [1:0] reg_rva_out_reg_data_30_25_sva_dfm_5_ftd_1;
  wire weight_port_read_out_data_0_1_sva_mx0_15;
  wire [14:0] weight_port_read_out_data_0_1_sva_mx0_14_0;
  wire rva_out_reg_data_and_130_ssc;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_1_3_2;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_1_1_0;
  wire weight_mem_run_3_for_5_and_158_ssc;
  wire weight_mem_run_3_for_5_and_159_ssc;
  wire weight_mem_run_3_for_5_and_160_ssc;
  wire weight_mem_run_3_for_5_and_161_ssc;
  wire weight_mem_run_3_for_5_and_164_ssc;
  wire weight_port_read_out_data_and_128_ssc;
  reg weight_port_read_out_data_0_1_sva_dfm_1_1_15;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_1_1_14_0;
  reg weight_port_read_out_data_0_1_sva_15;
  reg [14:0] weight_port_read_out_data_0_1_sva_14_0;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_2_3_2;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_2_1_0;
  reg weight_port_read_out_data_0_1_sva_dfm_4_15;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_4_14_0;
  wire rva_out_reg_data_and_89_ssc;
  reg [3:0] rva_out_reg_data_30_25_sva_dfm_6_5_2;
  reg [1:0] rva_out_reg_data_30_25_sva_dfm_6_1_0;
  wire [1:0] rva_out_reg_data_35_32_sva_dfm_6_mx1_3_2;
  wire [1:0] rva_out_reg_data_35_32_sva_dfm_6_mx1_1_0;
  wire rva_out_reg_data_and_26_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_2_cse;
  wire rva_out_reg_data_and_29_cse;
  wire input_mem_banks_read_read_data_and_cse;
  wire weight_port_read_out_data_and_125_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_cse;
  wire PECore_PushOutput_if_and_cse;
  wire rva_in_reg_rw_and_cse;
  wire PECore_RunMac_if_and_1_cse;
  wire PECore_RunMac_if_and_2_cse;
  wire input_mem_banks_read_1_read_data_and_cse;
  wire weight_mem_run_3_for_aelse_and_cse;
  wire data_in_tmp_operator_2_for_and_1_cse;
  wire data_in_tmp_operator_2_for_and_16_cse;
  wire PECore_RunMac_if_and_6_cse;
  wire weight_mem_run_3_for_aelse_and_5_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_52_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_58_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_64_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_69_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_74_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_79_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_85_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_90_cse;
  wire weight_read_addrs_and_4_cse;
  wire weight_write_data_data_and_cse;
  wire weight_mem_write_arbxbar_xbar_for_1_for_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse;
  wire PECore_RunFSM_switch_lp_and_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_15_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_22_cse;
  wire Arbiter_8U_Roundrobin_pick_and_85_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_64_cse;
  wire weight_write_data_data_and_16_cse;
  wire rva_in_reg_rw_and_4_cse;
  wire PECore_UpdateFSM_switch_lp_and_9_cse;
  wire state_and_cse;
  wire weight_port_read_out_data_and_131_cse;
  wire weight_read_addrs_and_15_cse;
  wire weight_read_addrs_and_16_cse;
  wire weight_port_read_out_data_and_134_cse;
  wire weight_port_read_out_data_and_150_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_374_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_378_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_382_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_387_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_389_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse;
  wire while_if_and_12_cse;
  wire weight_read_addrs_and_19_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse;
  wire rva_in_reg_rw_and_6_cse;
  wire input_mem_banks_read_read_data_and_9_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse;
  wire while_if_and_16_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_7_cse;
  wire while_if_and_6_cse;
  wire rva_out_reg_data_and_47_cse;
  wire weight_port_read_out_data_and_164_cse;
  wire input_read_req_valid_and_1_cse;
  wire weight_mem_banks_load_store_for_else_and_cse;
  wire weight_mem_banks_load_store_for_else_and_72_cse;
  wire weight_mem_banks_load_store_for_else_and_73_cse;
  wire weight_mem_banks_load_store_for_else_and_74_cse;
  wire weight_mem_banks_load_store_for_else_and_75_cse;
  wire rva_in_reg_rw_and_9_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_396_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_398_cse;
  wire weight_read_addrs_and_23_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_402_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_159_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_163_cse;
  wire input_mem_banks_read_read_data_and_18_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse;
  wire pe_manager_base_weight_and_5_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_11_cse;
  wire while_if_and_7_cse;
  wire rva_out_reg_data_and_68_cse;
  wire weight_port_read_out_data_and_166_cse;
  wire input_read_req_valid_and_2_cse;
  wire rva_in_reg_rw_and_5_cse;
  wire PECore_RunMac_if_and_3_cse;
  wire rva_in_reg_rw_and_12_cse;
  wire input_mem_banks_read_read_data_and_27_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_15_cse;
  wire while_if_and_8_cse;
  wire weight_port_read_out_data_and_168_cse;
  wire input_read_req_valid_and_3_cse;
  wire PECore_UpdateFSM_switch_lp_and_16_cse;
  wire PECore_RunMac_if_and_4_cse;
  wire rva_in_reg_rw_and_15_cse;
  wire input_mem_banks_read_read_data_and_36_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_19_cse;
  wire while_if_and_9_cse;
  wire input_read_req_valid_and_4_cse;
  wire PECore_UpdateFSM_switch_lp_and_18_cse;
  wire PECore_RunMac_if_and_5_cse;
  wire input_mem_banks_read_read_data_and_45_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_23_cse;
  wire rva_out_reg_data_and_128_cse;
  wire rva_out_reg_data_and_134_cse;
  wire input_read_req_valid_and_5_cse;
  wire rva_out_reg_data_and_146_cse;
  wire rva_out_reg_data_and_150_cse;
  wire PECore_RunMac_if_and_8_cse;
  wire rva_in_reg_rw_and_2_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_24_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_27_cse;
  wire rva_out_reg_data_and_166_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_28_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_31_cse;
  wire rva_out_reg_data_and_169_cse;
  wire rva_out_reg_data_and_172_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_33_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse;
  wire rva_out_reg_data_and_175_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_46_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_48_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_52_cse;
  wire weight_port_read_out_data_and_170_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_29_cse;
  wire accum_vector_data_and_16_cse;
  reg weight_port_read_out_data_0_1_sva_dfm_5_rsp_0;
  reg [14:0] weight_port_read_out_data_0_1_sva_dfm_5_rsp_1;
  reg [3:0] rva_out_reg_data_30_25_sva_dfm_7_rsp_0;
  reg [1:0] rva_out_reg_data_30_25_sva_dfm_7_rsp_1;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_3_rsp_0;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_3_rsp_1;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_6_rsp_0;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_6_rsp_1;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd;
  reg [14:0] reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd_1;
  reg [3:0] reg_rva_out_reg_data_30_25_sva_dfm_8_ftd;
  reg [1:0] reg_rva_out_reg_data_30_25_sva_dfm_8_ftd_1;
  reg [1:0] reg_rva_out_reg_data_35_32_sva_dfm_4_4_ftd;
  reg [1:0] reg_rva_out_reg_data_35_32_sva_dfm_4_4_ftd_1;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_5_3_2;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_5_1_0;
  reg [3:0] rva_out_reg_data_30_25_sva_dfm_9_5_2;
  reg [1:0] rva_out_reg_data_30_25_sva_dfm_9_1_0;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_6_rsp_0;
  reg [1:0] rva_out_reg_data_35_32_sva_dfm_4_6_rsp_1;
  wire [3:0] rva_out_reg_data_30_25_sva_dfm_7_5_2;
  wire [1:0] rva_out_reg_data_30_25_sva_dfm_7_1_0;
  reg [3:0] rva_out_reg_data_30_25_sva_dfm_6_5_2_1;
  reg [1:0] rva_out_reg_data_30_25_sva_dfm_6_1_0_1;
  wire and_dcpl_808;
  wire or_dcpl_752;
  wire or_dcpl_753;
  wire or_dcpl_761;
  wire or_dcpl_766;
  wire or_dcpl_774;
  wire or_dcpl_792;
  wire or_tmp_441;
  wire mux_tmp_376;
  wire and_1072_cse;
  wire and_1099_cse;
  wire or_1189_cse;
  wire and_1135_cse;
  wire and_1130_cse;
  wire xor_1_cse;
  wire and_1210_cse;
  wire or_1293_cse;
  wire nor_523_cse;
  wire nand_72_cse;
  wire nor_526_cse;
  wire nor_521_cse;
  wire nor_534_cse;
  wire nor_518_cse;
  wire nor_520_cse;
  wire and_1344_cse;
  wire or_666_cse;
  wire mux_403_cse;
  wire and_1441_cse;
  wire and_1227_cse;
  wire and_1437_cse;
  wire nor_500_cse;
  wire nor_508_cse;
  wire nand_83_cse;
  wire or_1284_cse;
  wire and_1141_cse;
  wire and_1156_cse;
  wire and_1165_cse;
  wire and_1201_cse;
  wire and_1294_cse;
  wire and_1357_cse;
  wire and_1372_cse;
  wire mux_402_cse;
  wire and_1266_cse;
  reg reg_rva_out_reg_data_15_9_sva_dfm_10_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_8_enexo;
  reg reg_rva_out_reg_data_255_240_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_239_224_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_223_208_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_207_192_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_191_176_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_175_160_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_159_144_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_143_128_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_127_112_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_111_96_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_95_80_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_5_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_4_5_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_5_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_5_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5_enexo;
  reg reg_accum_vector_data_6_35_0_sva_dfm_1_1_enexo;
  reg reg_accum_vector_data_5_35_0_sva_dfm_1_1_enexo;
  reg reg_accum_vector_data_4_35_0_sva_dfm_1_1_enexo;
  reg reg_accum_vector_data_3_35_0_sva_dfm_1_1_enexo;
  reg reg_accum_vector_data_2_35_0_sva_dfm_1_1_enexo;
  reg reg_accum_vector_data_1_35_0_sva_dfm_1_1_enexo;
  reg reg_accum_vector_data_0_35_0_sva_dfm_1_1_enexo;
  reg reg_accum_vector_data_7_35_0_sva_dfm_1_1_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000001;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000002;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000003;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000004;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000005;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000006;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000007;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000008;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000009;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000010;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000011;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000012;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000013;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000014;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000001;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000002;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000003;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000004;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000005;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000006;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000007;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000008;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000009;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000010;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000011;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000012;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000013;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000014;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2;
  reg reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1;
  reg reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  reg reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_addrs_lpi_1_dfm_1_1_enexo;
  reg reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_config_num_output_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  reg reg_rva_in_reg_data_sva_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_7_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_7_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_9_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_255_240_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_239_224_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_223_208_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_207_192_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_191_176_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_175_160_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_159_144_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_143_128_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_127_112_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_111_96_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_95_80_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_4_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_255_240_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_239_224_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_223_208_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_207_192_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_191_176_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_175_160_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_159_144_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_143_128_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_127_112_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_111_96_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_95_80_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_4_3_enexo;
  reg reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_2_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_255_240_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_239_224_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_223_208_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_207_192_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_191_176_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_175_160_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_159_144_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_143_128_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_127_112_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_111_96_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_95_80_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_4_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_6_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_255_240_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_239_224_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_223_208_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_207_192_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_191_176_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_175_160_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_159_144_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_143_128_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_127_112_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_111_96_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_95_80_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_79_64_sva_dfm_4_1_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_3;
  reg reg_rva_out_reg_data_23_17_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_4_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_1_3_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1;
  reg reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_62_48_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  reg reg_pe_manager_base_input_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_8_enexo;
  wire rva_out_reg_data_and_191_enex5;
  wire rva_out_reg_data_and_192_enex5;
  wire rva_out_reg_data_and_193_enex5;
  wire rva_out_reg_data_and_194_enex5;
  wire rva_out_reg_data_and_195_enex5;
  wire rva_out_reg_data_and_196_enex5;
  wire rva_out_reg_data_and_197_enex5;
  wire rva_out_reg_data_and_198_enex5;
  wire rva_out_reg_data_and_199_enex5;
  wire rva_out_reg_data_and_200_enex5;
  wire rva_out_reg_data_and_201_enex5;
  wire rva_out_reg_data_and_202_enex5;
  wire rva_out_reg_data_and_203_enex5;
  wire rva_out_reg_data_and_204_enex5;
  wire rva_out_reg_data_and_205_enex5;
  wire rva_out_reg_data_and_206_enex5;
  wire rva_out_reg_data_and_207_enex5;
  wire weight_port_read_out_data_and_172_enex5;
  wire input_mem_banks_read_read_data_and_57_enex5;
  wire input_mem_banks_read_read_data_and_58_enex5;
  wire weight_port_read_out_data_and_173_enex5;
  wire input_mem_banks_read_read_data_and_59_enex5;
  wire input_mem_banks_read_read_data_and_60_enex5;
  wire accum_vector_data_and_24_enex5;
  wire accum_vector_data_and_25_enex5;
  wire accum_vector_data_and_26_enex5;
  wire accum_vector_data_and_27_enex5;
  wire accum_vector_data_and_28_enex5;
  wire accum_vector_data_and_29_enex5;
  wire accum_vector_data_and_30_enex5;
  wire accum_vector_data_and_7_enex5;
  wire input_mem_banks_read_1_read_data_and_5_enex5;
  wire weight_port_read_out_data_and_enex5;
  wire weight_port_read_out_data_and_174_enex5;
  wire weight_port_read_out_data_and_175_enex5;
  wire weight_port_read_out_data_and_176_enex5;
  wire weight_port_read_out_data_and_177_enex5;
  wire weight_port_read_out_data_and_178_enex5;
  wire weight_port_read_out_data_and_179_enex5;
  wire weight_port_read_out_data_and_180_enex5;
  wire weight_port_read_out_data_and_181_enex5;
  wire weight_port_read_out_data_and_182_enex5;
  wire weight_port_read_out_data_and_183_enex5;
  wire weight_port_read_out_data_and_184_enex5;
  wire weight_port_read_out_data_and_185_enex5;
  wire weight_port_read_out_data_and_186_enex5;
  wire weight_port_read_out_data_and_187_enex5;
  wire weight_port_read_out_data_and_188_enex5;
  wire weight_port_read_out_data_and_189_enex5;
  wire weight_port_read_out_data_and_190_enex5;
  wire weight_port_read_out_data_and_191_enex5;
  wire weight_port_read_out_data_and_192_enex5;
  wire weight_port_read_out_data_and_193_enex5;
  wire weight_port_read_out_data_and_194_enex5;
  wire weight_port_read_out_data_and_195_enex5;
  wire weight_port_read_out_data_and_196_enex5;
  wire weight_port_read_out_data_and_197_enex5;
  wire weight_port_read_out_data_and_198_enex5;
  wire weight_port_read_out_data_and_199_enex5;
  wire weight_port_read_out_data_and_200_enex5;
  wire weight_port_read_out_data_and_201_enex5;
  wire weight_port_read_out_data_and_202_enex5;
  wire weight_port_read_out_data_and_203_enex5;
  wire weight_port_read_out_data_and_31_enex5;
  wire input_mem_banks_read_1_read_data_and_1_enex5;
  wire weight_read_addrs_and_2_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5;
  wire weight_write_data_data_and_48_enex5;
  wire weight_write_data_data_and_49_enex5;
  wire weight_write_data_data_and_50_enex5;
  wire weight_write_data_data_and_51_enex5;
  wire weight_write_data_data_and_52_enex5;
  wire weight_write_data_data_and_53_enex5;
  wire weight_write_data_data_and_54_enex5;
  wire weight_write_data_data_and_55_enex5;
  wire weight_write_data_data_and_56_enex5;
  wire weight_write_data_data_and_57_enex5;
  wire weight_write_data_data_and_58_enex5;
  wire weight_write_data_data_and_59_enex5;
  wire weight_write_data_data_and_60_enex5;
  wire weight_write_data_data_and_61_enex5;
  wire weight_write_data_data_and_62_enex5;
  wire weight_write_data_data_and_63_enex5;
  wire weight_write_addrs_and_enex5;
  wire weight_write_data_data_and_64_enex5;
  wire weight_write_data_data_and_65_enex5;
  wire weight_write_data_data_and_66_enex5;
  wire weight_write_data_data_and_67_enex5;
  wire weight_write_data_data_and_68_enex5;
  wire weight_write_data_data_and_69_enex5;
  wire weight_write_data_data_and_70_enex5;
  wire weight_write_data_data_and_71_enex5;
  wire weight_write_data_data_and_72_enex5;
  wire weight_write_data_data_and_73_enex5;
  wire weight_write_data_data_and_74_enex5;
  wire weight_write_data_data_and_75_enex5;
  wire weight_write_data_data_and_76_enex5;
  wire weight_write_data_data_and_77_enex5;
  wire weight_write_data_data_and_78_enex5;
  wire weight_write_data_data_and_79_enex5;
  wire weight_write_addrs_and_3_enex5;
  wire weight_read_addrs_and_enex5;
  wire pe_config_UpdateManagerCounter_if_if_and_enex5;
  wire weight_read_addrs_and_27_enex5;
  wire PEManager_15U_PEManagerWrite_and_enex5;
  wire input_mem_banks_read_read_data_and_61_enex5;
  wire input_mem_banks_read_read_data_and_62_enex5;
  wire input_mem_banks_read_read_data_and_63_enex5;
  wire input_mem_banks_read_read_data_and_64_enex5;
  wire input_mem_banks_read_1_read_data_and_2_enex5;
  wire rva_out_reg_data_and_208_enex5;
  wire rva_out_reg_data_and_209_enex5;
  wire rva_out_reg_data_and_210_enex5;
  wire weight_port_read_out_data_and_204_enex5;
  wire rva_out_reg_data_and_211_enex5;
  wire rva_out_reg_data_and_212_enex5;
  wire rva_out_reg_data_and_213_enex5;
  wire rva_out_reg_data_and_214_enex5;
  wire rva_out_reg_data_and_215_enex5;
  wire rva_out_reg_data_and_216_enex5;
  wire rva_out_reg_data_and_217_enex5;
  wire rva_out_reg_data_and_218_enex5;
  wire rva_out_reg_data_and_219_enex5;
  wire rva_out_reg_data_and_220_enex5;
  wire rva_out_reg_data_and_221_enex5;
  wire rva_out_reg_data_and_222_enex5;
  wire rva_out_reg_data_and_223_enex5;
  wire rva_out_reg_data_and_224_enex5;
  wire rva_out_reg_data_and_225_enex5;
  wire input_mem_banks_read_read_data_and_65_enex5;
  wire input_mem_banks_read_read_data_and_66_enex5;
  wire input_mem_banks_read_read_data_and_67_enex5;
  wire input_mem_banks_read_read_data_and_68_enex5;
  wire input_mem_banks_read_1_read_data_and_3_enex5;
  wire rva_out_reg_data_and_226_enex5;
  wire rva_out_reg_data_and_227_enex5;
  wire weight_port_read_out_data_and_205_enex5;
  wire rva_out_reg_data_and_228_enex5;
  wire rva_out_reg_data_and_229_enex5;
  wire rva_out_reg_data_and_230_enex5;
  wire rva_out_reg_data_and_231_enex5;
  wire rva_out_reg_data_and_232_enex5;
  wire rva_out_reg_data_and_233_enex5;
  wire rva_out_reg_data_and_234_enex5;
  wire rva_out_reg_data_and_235_enex5;
  wire rva_out_reg_data_and_236_enex5;
  wire rva_out_reg_data_and_237_enex5;
  wire rva_out_reg_data_and_238_enex5;
  wire rva_out_reg_data_and_239_enex5;
  wire rva_out_reg_data_and_240_enex5;
  wire rva_out_reg_data_and_241_enex5;
  wire rva_out_reg_data_and_242_enex5;
  wire weight_mem_write_arbxbar_xbar_for_empty_and_3_enex5;
  wire input_mem_banks_read_read_data_and_69_enex5;
  wire input_mem_banks_read_read_data_and_70_enex5;
  wire input_mem_banks_read_read_data_and_71_enex5;
  wire input_mem_banks_read_read_data_and_72_enex5;
  wire rva_out_reg_data_and_243_enex5;
  wire rva_out_reg_data_and_244_enex5;
  wire weight_port_read_out_data_and_206_enex5;
  wire weight_port_read_out_data_and_207_enex5;
  wire rva_out_reg_data_and_245_enex5;
  wire rva_out_reg_data_and_246_enex5;
  wire rva_out_reg_data_and_247_enex5;
  wire rva_out_reg_data_and_248_enex5;
  wire rva_out_reg_data_and_249_enex5;
  wire rva_out_reg_data_and_250_enex5;
  wire rva_out_reg_data_and_251_enex5;
  wire rva_out_reg_data_and_252_enex5;
  wire rva_out_reg_data_and_253_enex5;
  wire rva_out_reg_data_and_254_enex5;
  wire rva_out_reg_data_and_255_enex5;
  wire rva_out_reg_data_and_256_enex5;
  wire rva_out_reg_data_and_257_enex5;
  wire rva_out_reg_data_and_258_enex5;
  wire rva_out_reg_data_and_259_enex5;
  wire input_mem_banks_read_read_data_and_73_enex5;
  wire input_mem_banks_read_read_data_and_74_enex5;
  wire input_mem_banks_read_read_data_and_75_enex5;
  wire input_mem_banks_read_read_data_and_76_enex5;
  wire rva_out_reg_data_and_260_enex5;
  wire rva_out_reg_data_and_261_enex5;
  wire rva_out_reg_data_and_262_enex5;
  wire weight_port_read_out_data_and_208_enex5;
  wire rva_out_reg_data_and_263_enex5;
  wire rva_out_reg_data_and_264_enex5;
  wire rva_out_reg_data_and_265_enex5;
  wire rva_out_reg_data_and_266_enex5;
  wire rva_out_reg_data_and_267_enex5;
  wire rva_out_reg_data_and_268_enex5;
  wire rva_out_reg_data_and_269_enex5;
  wire rva_out_reg_data_and_270_enex5;
  wire rva_out_reg_data_and_271_enex5;
  wire rva_out_reg_data_and_272_enex5;
  wire rva_out_reg_data_and_273_enex5;
  wire rva_out_reg_data_and_274_enex5;
  wire rva_out_reg_data_and_275_enex5;
  wire rva_out_reg_data_and_276_enex5;
  wire rva_out_reg_data_and_277_enex5;
  wire input_mem_banks_read_read_data_and_77_enex5;
  wire input_mem_banks_read_read_data_and_78_enex5;
  wire input_mem_banks_read_read_data_and_79_enex5;
  wire input_mem_banks_read_read_data_and_80_enex5;
  wire rva_out_reg_data_and_278_enex5;
  wire rva_out_reg_data_and_279_enex5;
  wire rva_out_reg_data_and_280_enex5;
  wire rva_out_reg_data_and_281_enex5;
  wire rva_out_reg_data_and_282_enex5;
  wire rva_out_reg_data_and_283_enex5;
  wire input_mem_banks_read_read_data_and_55_enex5;
  wire rva_out_reg_data_and_284_enex5;
  wire rva_out_reg_data_and_285_enex5;
  wire rva_out_reg_data_and_286_enex5;
  wire rva_out_reg_data_and_287_enex5;
  wire rva_out_reg_data_and_288_enex5;
  wire input_mem_banks_read_read_data_and_56_enex5;
  wire rva_out_reg_data_and_289_enex5;
  wire rva_out_reg_data_and_290_enex5;
  wire rva_out_reg_data_and_291_enex5;
  wire rva_out_reg_data_and_292_enex5;
  wire rva_out_reg_data_and_293_enex5;
  wire rva_out_reg_data_and_182_enex5;
  wire rva_out_reg_data_and_294_enex5;
  wire rva_out_reg_data_and_295_enex5;
  wire rva_out_reg_data_and_296_enex5;
  wire rva_out_reg_data_and_297_enex5;
  wire weight_port_read_out_data_and_209_enex5;
  wire rva_out_reg_data_and_298_enex5;
  wire rva_out_reg_data_and_299_enex5;
  wire rva_out_reg_data_and_300_enex5;
  wire weight_port_read_out_data_and_210_enex5;
  wire rva_out_reg_data_and_301_enex5;
  wire weight_port_read_out_data_and_211_enex5;
  wire rva_out_reg_data_and_302_enex5;
  wire rva_out_reg_data_and_303_enex5;
  wire and_1120_tmp;
  wire data_in_tmp_operator_2_for_and_tmp;
  wire data_in_tmp_operator_2_for_and_31_tmp;
  wire rva_in_reg_data_and_tmp;
  wire input_mem_banks_read_1_read_data_and_4_tmp;
  wire weight_port_read_out_data_and_127_tmp;
  wire input_mem_banks_read_read_data_and_54_tmp;
  wire pe_manager_base_input_and_tmp;
  wire rva_in_reg_rw_and_3_cse;
  wire and_1065_itm;
  wire and_756_itm;
  wire while_mux_1457_cse_1;
  wire while_mux_1429_cse_1;
  wire and_768_cse;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27;
  wire mux_70_nl;
  wire and_540_nl;
  wire nor_18_nl;
  wire mux_73_nl;
  wire mux_72_nl;
  wire or_697_nl;
  wire mux_71_nl;
  wire and_543_nl;
  wire and_988_nl;
  wire mux_76_nl;
  wire or_700_nl;
  wire mux_75_nl;
  wire nand_nl;
  wire mux_82_nl;
  wire mux_81_nl;
  wire mux_80_nl;
  wire or_706_nl;
  wire mux_79_nl;
  wire mux_78_nl;
  wire or_705_nl;
  wire or_704_nl;
  wire or_703_nl;
  wire mux_85_nl;
  wire mux_84_nl;
  wire or_710_nl;
  wire or_709_nl;
  wire mux_88_nl;
  wire mux_87_nl;
  wire or_718_nl;
  wire or_1149_nl;
  wire mux_91_nl;
  wire mux_90_nl;
  wire or_722_nl;
  wire or_1150_nl;
  wire mux_94_nl;
  wire or_726_nl;
  wire mux_93_nl;
  wire nand_3_nl;
  wire mux_98_nl;
  wire or_735_nl;
  wire mux_97_nl;
  wire nand_4_nl;
  wire mux_101_nl;
  wire mux_100_nl;
  wire or_739_nl;
  wire or_1151_nl;
  wire mux_114_nl;
  wire mux_113_nl;
  wire mux_112_nl;
  wire mux_111_nl;
  wire mux_110_nl;
  wire mux_467_nl;
  wire and_767_nl;
  wire mux_106_nl;
  wire mux_349_nl;
  wire mux_109_nl;
  wire mux_108_nl;
  wire mux_107_nl;
  wire mux_468_nl;
  wire mux_469_nl;
  wire or_140_nl;
  wire or_139_nl;
  wire or_138_nl;
  wire or_137_nl;
  wire PECore_UpdateFSM_switch_lp_not_25_nl;
  wire PECore_UpdateFSM_switch_lp_not_26_nl;
  wire PECore_UpdateFSM_switch_lp_not_27_nl;
  wire PECore_UpdateFSM_switch_lp_not_28_nl;
  wire PECore_UpdateFSM_switch_lp_not_29_nl;
  wire PECore_UpdateFSM_switch_lp_not_30_nl;
  wire PECore_UpdateFSM_switch_lp_not_19_nl;
  wire[35:0] PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_nl;
  wire[35:0] ProductSum_for_acc_40_nl;
  wire[37:0] nl_ProductSum_for_acc_40_nl;
  wire[35:0] ProductSum_for_acc_41_nl;
  wire[37:0] nl_ProductSum_for_acc_41_nl;
  wire[35:0] ProductSum_for_acc_42_nl;
  wire[37:0] nl_ProductSum_for_acc_42_nl;
  wire[34:0] ProductSum_for_acc_43_nl;
  wire[35:0] nl_ProductSum_for_acc_43_nl;
  wire PECore_UpdateFSM_switch_lp_not_31_nl;
  wire[35:0] PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_1_nl;
  wire[35:0] ProductSum_for_acc_32_nl;
  wire[37:0] nl_ProductSum_for_acc_32_nl;
  wire[35:0] ProductSum_for_acc_33_nl;
  wire[37:0] nl_ProductSum_for_acc_33_nl;
  wire[35:0] ProductSum_for_acc_34_nl;
  wire[37:0] nl_ProductSum_for_acc_34_nl;
  wire[34:0] ProductSum_for_acc_35_nl;
  wire[35:0] nl_ProductSum_for_acc_35_nl;
  wire PECore_UpdateFSM_switch_lp_not_32_nl;
  wire[35:0] PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_2_nl;
  wire[35:0] ProductSum_for_acc_24_nl;
  wire[37:0] nl_ProductSum_for_acc_24_nl;
  wire[35:0] ProductSum_for_acc_25_nl;
  wire[37:0] nl_ProductSum_for_acc_25_nl;
  wire[35:0] ProductSum_for_acc_26_nl;
  wire[37:0] nl_ProductSum_for_acc_26_nl;
  wire[34:0] ProductSum_for_acc_27_nl;
  wire[35:0] nl_ProductSum_for_acc_27_nl;
  wire PECore_UpdateFSM_switch_lp_not_33_nl;
  wire[35:0] PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_3_nl;
  wire[35:0] ProductSum_for_acc_20_nl;
  wire[37:0] nl_ProductSum_for_acc_20_nl;
  wire[35:0] ProductSum_for_acc_21_nl;
  wire[37:0] nl_ProductSum_for_acc_21_nl;
  wire[35:0] ProductSum_for_acc_22_nl;
  wire[37:0] nl_ProductSum_for_acc_22_nl;
  wire[34:0] ProductSum_for_acc_23_nl;
  wire[35:0] nl_ProductSum_for_acc_23_nl;
  wire PECore_UpdateFSM_switch_lp_not_34_nl;
  wire[35:0] PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_4_nl;
  wire[35:0] ProductSum_for_acc_28_nl;
  wire[37:0] nl_ProductSum_for_acc_28_nl;
  wire[35:0] ProductSum_for_acc_29_nl;
  wire[37:0] nl_ProductSum_for_acc_29_nl;
  wire[35:0] ProductSum_for_acc_30_nl;
  wire[37:0] nl_ProductSum_for_acc_30_nl;
  wire[34:0] ProductSum_for_acc_31_nl;
  wire[35:0] nl_ProductSum_for_acc_31_nl;
  wire PECore_UpdateFSM_switch_lp_not_35_nl;
  wire[35:0] PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_5_nl;
  wire[35:0] ProductSum_for_acc_36_nl;
  wire[37:0] nl_ProductSum_for_acc_36_nl;
  wire[35:0] ProductSum_for_acc_37_nl;
  wire[37:0] nl_ProductSum_for_acc_37_nl;
  wire[35:0] ProductSum_for_acc_38_nl;
  wire[37:0] nl_ProductSum_for_acc_38_nl;
  wire[34:0] ProductSum_for_acc_39_nl;
  wire[35:0] nl_ProductSum_for_acc_39_nl;
  wire PECore_UpdateFSM_switch_lp_not_36_nl;
  wire[35:0] PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_6_nl;
  wire[35:0] ProductSum_for_acc_44_nl;
  wire[37:0] nl_ProductSum_for_acc_44_nl;
  wire[35:0] ProductSum_for_acc_45_nl;
  wire[37:0] nl_ProductSum_for_acc_45_nl;
  wire[35:0] ProductSum_for_acc_46_nl;
  wire[37:0] nl_ProductSum_for_acc_46_nl;
  wire[34:0] ProductSum_for_acc_47_nl;
  wire[35:0] nl_ProductSum_for_acc_47_nl;
  wire PECore_UpdateFSM_switch_lp_not_21_nl;
  wire[35:0] PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_7_nl;
  wire[35:0] ProductSum_for_acc_nl;
  wire[37:0] nl_ProductSum_for_acc_nl;
  wire[35:0] ProductSum_for_acc_48_nl;
  wire[37:0] nl_ProductSum_for_acc_48_nl;
  wire[35:0] ProductSum_for_acc_49_nl;
  wire[37:0] nl_ProductSum_for_acc_49_nl;
  wire[34:0] ProductSum_for_acc_50_nl;
  wire[35:0] nl_ProductSum_for_acc_50_nl;
  wire PECore_UpdateFSM_switch_lp_not_10_nl;
  wire weight_mem_run_3_for_5_and_166_nl;
  wire weight_mem_run_3_for_5_and_167_nl;
  wire weight_mem_run_3_for_5_and_168_nl;
  wire weight_mem_run_3_for_5_and_169_nl;
  wire weight_mem_run_3_for_5_and_170_nl;
  wire weight_mem_run_3_for_5_and_172_nl;
  wire mux_354_nl;
  wire or_1188_nl;
  wire weight_mem_run_3_for_5_and_174_nl;
  wire weight_mem_run_3_for_5_and_175_nl;
  wire weight_mem_run_3_for_5_and_176_nl;
  wire weight_mem_run_3_for_5_and_177_nl;
  wire weight_mem_run_3_for_5_and_179_nl;
  wire weight_mem_run_3_for_5_and_180_nl;
  wire mux_355_nl;
  wire or_1190_nl;
  wire[15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl;
  wire[15:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_1_nl;
  wire mux_357_nl;
  wire mux_356_nl;
  wire mux_373_nl;
  wire mux_372_nl;
  wire mux_376_nl;
  wire nor_510_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_48_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl;
  wire mux_5_nl;
  wire mux_4_nl;
  wire and_64_nl;
  wire and_766_nl;
  wire or_13_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_80_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_138_nl;
  wire mux_6_nl;
  wire nor_328_nl;
  wire mux_7_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_80_nl;
  wire mux_378_nl;
  wire mux_377_nl;
  wire nor_511_nl;
  wire nor_512_nl;
  wire[10:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl;
  wire[3:0] PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl;
  wire and_622_nl;
  wire[3:0] operator_4_false_acc_nl;
  wire[4:0] nl_operator_4_false_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_7_nl;
  wire mux_379_nl;
  wire mux_380_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_and_1_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_mux1h_16_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_nor_8_nl;
  wire PECore_UpdateFSM_switch_lp_not_11_nl;
  wire mux_390_nl;
  wire nor_525_nl;
  wire mux_393_nl;
  wire or_1318_nl;
  wire mux_392_nl;
  wire mux_391_nl;
  wire mux_396_nl;
  wire mux_395_nl;
  wire mux_394_nl;
  wire or_1326_nl;
  wire or_1325_nl;
  wire or_1324_nl;
  wire mux_36_nl;
  wire mux_3_nl;
  wire mux_2_nl;
  wire nor_273_nl;
  wire or_8_nl;
  wire mux_399_nl;
  wire or_1335_nl;
  wire or_1333_nl;
  wire mux_398_nl;
  wire mux_397_nl;
  wire and_1442_nl;
  wire and_1443_nl;
  wire and_1444_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_nl;
  wire mux_37_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_136_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_215_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_18_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_204_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_28_nl;
  wire mux_41_nl;
  wire mux_40_nl;
  wire or_189_nl;
  wire mux_38_nl;
  wire or_182_nl;
  wire or_180_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_27_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_234_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_249_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_174_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_189_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_204_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_219_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_235_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_250_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_175_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_190_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_205_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_220_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_236_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_251_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_176_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_191_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_206_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_221_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_237_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_252_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_177_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_192_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_207_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_222_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_238_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_253_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_178_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_193_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_208_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_223_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_239_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_254_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_179_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_194_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_209_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_224_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_240_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_255_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_180_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_195_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_210_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_225_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_241_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_181_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_196_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_211_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_226_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_242_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_257_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_182_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_197_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_212_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_227_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_243_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_183_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_198_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_213_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_228_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_244_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_259_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_184_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_199_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_214_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_229_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_245_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_260_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_185_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_200_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_215_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_230_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_246_nl;
  wire mux_43_nl;
  wire mux_42_nl;
  wire nor_291_nl;
  wire[15:0] mux1h_2_nl;
  wire not_2436_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_201_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_231_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_247_nl;
  wire[15:0] mux1h_3_nl;
  wire not_2438_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_202_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_232_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_248_nl;
  wire[15:0] mux1h_4_nl;
  wire not_2440_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_203_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_233_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_140_nl;
  wire[15:0] mux_348_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_or_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_mux1h_89_nl;
  wire and_669_nl;
  wire and_670_nl;
  wire and_672_nl;
  wire and_675_nl;
  wire and_678_nl;
  wire and_668_nl;
  wire mux_340_nl;
  wire and_1061_nl;
  wire nor_471_nl;
  wire nand_67_nl;
  wire mux_49_nl;
  wire mux_48_nl;
  wire or_206_nl;
  wire mux_47_nl;
  wire or_205_nl;
  wire or_200_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_135_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_134_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_132_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_nl;
  wire mux_50_nl;
  wire mux_53_nl;
  wire mux_52_nl;
  wire nor_339_nl;
  wire[7:0] input_mem_banks_read_1_for_mux_nl;
  wire and_1062_nl;
  wire[14:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl;
  wire or_834_nl;
  wire mux_54_nl;
  wire or_160_nl;
  wire mux_55_nl;
  wire mux_61_nl;
  wire mux_60_nl;
  wire or_671_nl;
  wire mux_59_nl;
  wire mux_401_nl;
  wire mux_400_nl;
  wire or_1369_nl;
  wire or_1368_nl;
  wire or_1367_nl;
  wire or_1366_nl;
  wire or_1365_nl;
  wire mux_404_nl;
  wire weight_port_read_out_data_mux_67_nl;
  wire and_688_nl;
  wire nor_463_nl;
  wire mux_62_nl;
  wire mux_66_nl;
  wire mux_65_nl;
  wire mux_64_nl;
  wire mux_63_nl;
  wire and_762_nl;
  wire or_674_nl;
  wire mux_67_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_6_nl;
  wire PECore_PushAxiRsp_if_else_mux_27_nl;
  wire rva_out_reg_data_mux_34_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_21_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl;
  wire PECore_PushAxiRsp_if_else_mux_28_nl;
  wire rva_out_reg_data_mux_35_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_22_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_mux_18_nl;
  wire PECore_PushAxiRsp_if_else_mux_29_nl;
  wire rva_out_reg_data_mux_36_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_23_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl;
  wire[6:0] PECore_DecodeAxiRead_switch_lp_mux_19_nl;
  wire PECore_PushAxiRsp_if_else_mux_30_nl;
  wire rva_out_reg_data_mux_38_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_24_nl;
  wire[3:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl;
  wire[3:0] PECore_DecodeAxiRead_switch_lp_mux_20_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl;
  wire[1:0] PECore_DecodeAxiRead_switch_lp_mux_25_nl;
  wire PECore_PushAxiRsp_if_else_mux_31_nl;
  wire rva_out_reg_data_mux_37_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl;
  wire PECore_RunScale_and_14_nl;
  wire PECore_RunScale_and_15_nl;
  wire PECore_RunScale_and_12_nl;
  wire PECore_RunScale_and_13_nl;
  wire PECore_RunScale_and_10_nl;
  wire PECore_RunScale_and_11_nl;
  wire PECore_RunScale_and_8_nl;
  wire PECore_RunScale_and_9_nl;
  wire PECore_RunScale_and_6_nl;
  wire PECore_RunScale_and_7_nl;
  wire PECore_RunScale_and_4_nl;
  wire PECore_RunScale_and_5_nl;
  wire PECore_RunScale_and_2_nl;
  wire PECore_RunScale_and_3_nl;
  wire PECore_RunMac_or_nl;
  wire PECore_RunScale_and_nl;
  wire PECore_RunScale_and_1_nl;
  wire[15:0] mux1h_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_nl;
  wire not_2443_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_69_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_73_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_77_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_81_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_85_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_95_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_98_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_99_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_103_nl;
  wire[14:0] PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_nl;
  wire[14:0] nl_operator_15_false_acc_nl;
  wire[14:0] PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[12:0] operator_15_false_acc_1_nl;
  wire[13:0] nl_operator_15_false_acc_1_nl;
  wire[14:0] PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_2_nl;
  wire[14:0] nl_operator_15_false_acc_2_nl;
  wire[14:0] PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl;
  wire and_665_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl;
  wire and_658_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl;
  wire and_651_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl;
  wire and_644_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl;
  wire and_637_nl;
  wire[7:0] pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl;
  wire[7:0] operator_8_false_acc_nl;
  wire[8:0] nl_operator_8_false_acc_nl;
  wire pe_config_UpdateInputCounter_not_nl;
  wire pe_config_input_counter_nand_nl;
  wire[7:0] pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl;
  wire[7:0] operator_8_false_1_acc_nl;
  wire[8:0] nl_operator_8_false_1_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_9_nl;
  wire pe_config_output_counter_nand_nl;
  wire while_and_164_nl;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl;
  wire while_if_or_nl;
  wire while_if_and_4_nl;
  wire[15:0] mux1h_5_nl;
  wire not_2445_nl;
  wire[15:0] mux1h_6_nl;
  wire and_1053_nl;
  wire not_2447_nl;
  wire PECore_PushAxiRsp_mux_27_nl;
  wire[15:0] while_if_while_if_and_24_nl;
  wire[15:0] while_if_while_if_and_25_nl;
  wire[15:0] while_if_while_if_and_26_nl;
  wire[15:0] while_if_while_if_and_27_nl;
  wire[15:0] while_if_while_if_and_28_nl;
  wire[15:0] while_if_while_if_and_29_nl;
  wire[15:0] while_if_while_if_and_30_nl;
  wire[15:0] while_if_while_if_and_31_nl;
  wire[15:0] while_if_while_if_and_32_nl;
  wire[15:0] while_if_while_if_and_33_nl;
  wire[15:0] while_if_while_if_and_34_nl;
  wire[15:0] while_if_while_if_and_35_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_nl;
  wire weight_mem_banks_load_store_1_for_else_else_or_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_4_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_6_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_8_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_146_nl;
  wire mux_145_nl;
  wire mux_144_nl;
  wire or_887_nl;
  wire or_884_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_182_nl;
  wire mux_181_nl;
  wire mux_180_nl;
  wire or_934_nl;
  wire or_929_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl;
  wire and_707_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl;
  wire and_718_nl;
  wire mux_206_nl;
  wire nor_464_nl;
  wire nor_465_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_24_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl;
  wire and_732_nl;
  wire mux_240_nl;
  wire mux_239_nl;
  wire or_1010_nl;
  wire or_1009_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_286_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl;
  wire and_749_nl;
  wire mux_294_nl;
  wire nor_466_nl;
  wire nor_467_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_46_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_47_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_337_nl;
  wire mux_336_nl;
  wire or_1141_nl;
  wire mux_334_nl;
  wire or_1129_nl;
  wire PECore_UpdateFSM_switch_lp_mux1h_15_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl;
  wire PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl;
  wire PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_69_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_111_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_144_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_127_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_159_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_110_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_145_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_126_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_160_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_109_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_146_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_125_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_161_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_108_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_147_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_124_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_162_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_100_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_148_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_116_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_163_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_107_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_149_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_123_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_164_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_101_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_150_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_117_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_165_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_106_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_151_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_122_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_166_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_102_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_152_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_118_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_167_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_105_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_153_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_121_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_168_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_103_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_154_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_119_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_169_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_104_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_155_nl;
  wire[15:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_120_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_170_nl;
  wire[7:0] PEManager_15U_GetInputAddr_acc_nl;
  wire[8:0] nl_PEManager_15U_GetInputAddr_acc_nl;
  wire PECore_PushAxiRsp_mux_24_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_583_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_584_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_585_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_586_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_587_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_588_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_589_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_590_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_591_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_592_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_593_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_594_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_601_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_603_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_606_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_611_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_619_nl;
  wire mux_12_nl;
  wire mux_11_nl;
  wire mux_10_nl;
  wire and_753_nl;
  wire mux_45_nl;
  wire nand_29_nl;
  wire or_203_nl;
  wire or_202_nl;
  wire and_759_nl;
  wire mux_74_nl;
  wire or_698_nl;
  wire mux_77_nl;
  wire or_702_nl;
  wire mux_83_nl;
  wire or_708_nl;
  wire mux_86_nl;
  wire or_713_nl;
  wire mux_89_nl;
  wire or_721_nl;
  wire mux_92_nl;
  wire or_724_nl;
  wire mux_95_nl;
  wire or_732_nl;
  wire mux_96_nl;
  wire or_728_nl;
  wire mux_99_nl;
  wire or_738_nl;
  wire mux_125_nl;
  wire mux_124_nl;
  wire or_843_nl;
  wire or_841_nl;
  wire mux_128_nl;
  wire mux_127_nl;
  wire or_855_nl;
  wire or_849_nl;
  wire mux_135_nl;
  wire mux_134_nl;
  wire mux_133_nl;
  wire or_873_nl;
  wire or_871_nl;
  wire mux_132_nl;
  wire mux_131_nl;
  wire or_870_nl;
  wire or_868_nl;
  wire mux_130_nl;
  wire or_867_nl;
  wire or_861_nl;
  wire mux_143_nl;
  wire mux_142_nl;
  wire mux_141_nl;
  wire mux_140_nl;
  wire nor_384_nl;
  wire nor_385_nl;
  wire nor_386_nl;
  wire nor_387_nl;
  wire mux_139_nl;
  wire mux_138_nl;
  wire mux_137_nl;
  wire nor_388_nl;
  wire nor_389_nl;
  wire nor_390_nl;
  wire nor_391_nl;
  wire mux_148_nl;
  wire mux_147_nl;
  wire or_891_nl;
  wire or_889_nl;
  wire mux_151_nl;
  wire mux_150_nl;
  wire nand_6_nl;
  wire mux_154_nl;
  wire mux_153_nl;
  wire nand_7_nl;
  wire mux_157_nl;
  wire mux_156_nl;
  wire or_893_nl;
  wire or_892_nl;
  wire mux_161_nl;
  wire mux_160_nl;
  wire mux_159_nl;
  wire or_898_nl;
  wire or_897_nl;
  wire or_896_nl;
  wire mux_165_nl;
  wire mux_164_nl;
  wire mux_163_nl;
  wire or_905_nl;
  wire or_904_nl;
  wire mux_171_nl;
  wire mux_170_nl;
  wire mux_169_nl;
  wire or_912_nl;
  wire or_911_nl;
  wire mux_168_nl;
  wire mux_167_nl;
  wire or_910_nl;
  wire or_909_nl;
  wire mux_166_nl;
  wire or_908_nl;
  wire or_901_nl;
  wire mux_179_nl;
  wire mux_178_nl;
  wire mux_177_nl;
  wire mux_176_nl;
  wire nor_392_nl;
  wire nor_393_nl;
  wire nor_394_nl;
  wire nor_395_nl;
  wire mux_175_nl;
  wire mux_174_nl;
  wire mux_173_nl;
  wire nor_396_nl;
  wire nor_397_nl;
  wire nor_398_nl;
  wire nor_399_nl;
  wire mux_183_nl;
  wire while_mux_1482_nl;
  wire while_mux_1463_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_595_nl;
  wire mux_186_nl;
  wire mux_185_nl;
  wire mux_184_nl;
  wire nor_402_nl;
  wire nor_403_nl;
  wire or_943_nl;
  wire or_942_nl;
  wire mux_191_nl;
  wire mux_190_nl;
  wire nand_8_nl;
  wire or_941_nl;
  wire mux_199_nl;
  wire mux_198_nl;
  wire mux_197_nl;
  wire mux_196_nl;
  wire mux_195_nl;
  wire mux_194_nl;
  wire or_947_nl;
  wire mux_204_nl;
  wire nor_410_nl;
  wire mux_203_nl;
  wire or_956_nl;
  wire mux_202_nl;
  wire or_955_nl;
  wire nor_411_nl;
  wire mux_201_nl;
  wire or_952_nl;
  wire mux_200_nl;
  wire or_951_nl;
  wire mux_205_nl;
  wire nor_412_nl;
  wire nor_413_nl;
  wire mux_207_nl;
  wire while_mux_1446_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_610_nl;
  wire mux_210_nl;
  wire or_975_nl;
  wire nand_12_nl;
  wire mux_214_nl;
  wire mux_213_nl;
  wire mux_212_nl;
  wire or_974_nl;
  wire or_972_nl;
  wire mux_209_nl;
  wire mux_208_nl;
  wire or_971_nl;
  wire or_969_nl;
  wire mux_218_nl;
  wire mux_217_nl;
  wire mux_216_nl;
  wire nor_417_nl;
  wire nor_418_nl;
  wire mux_219_nl;
  wire or_986_nl;
  wire or_985_nl;
  wire or_983_nl;
  wire mux_224_nl;
  wire or_994_nl;
  wire mux_229_nl;
  wire mux_228_nl;
  wire nor_425_nl;
  wire mux_227_nl;
  wire mux_226_nl;
  wire nor_426_nl;
  wire nor_427_nl;
  wire mux_223_nl;
  wire nor_428_nl;
  wire mux_222_nl;
  wire or_992_nl;
  wire mux_221_nl;
  wire nor_429_nl;
  wire nor_430_nl;
  wire mux_232_nl;
  wire or_1006_nl;
  wire nand_16_nl;
  wire mux_236_nl;
  wire mux_235_nl;
  wire mux_234_nl;
  wire or_1005_nl;
  wire or_1003_nl;
  wire mux_231_nl;
  wire mux_230_nl;
  wire or_1002_nl;
  wire or_1000_nl;
  wire or_1011_nl;
  wire mux_246_nl;
  wire mux_245_nl;
  wire mux_244_nl;
  wire or_1016_nl;
  wire mux_243_nl;
  wire or_1015_nl;
  wire or_1013_nl;
  wire mux_249_nl;
  wire mux_248_nl;
  wire nand_17_nl;
  wire mux_256_nl;
  wire or_1023_nl;
  wire mux_255_nl;
  wire mux_254_nl;
  wire mux_253_nl;
  wire mux_252_nl;
  wire nand_18_nl;
  wire mux_251_nl;
  wire or_1019_nl;
  wire mux_258_nl;
  wire or_1025_nl;
  wire or_1024_nl;
  wire or_1035_nl;
  wire mux_261_nl;
  wire or_1032_nl;
  wire or_1037_nl;
  wire mux_263_nl;
  wire or_1036_nl;
  wire or_1030_nl;
  wire mux_265_nl;
  wire mux_268_nl;
  wire or_1040_nl;
  wire mux_267_nl;
  wire or_1039_nl;
  wire or_1038_nl;
  wire mux_275_nl;
  wire mux_274_nl;
  wire mux_273_nl;
  wire mux_272_nl;
  wire or_1051_nl;
  wire mux_271_nl;
  wire mux_270_nl;
  wire or_1048_nl;
  wire or_1047_nl;
  wire mux_269_nl;
  wire or_1046_nl;
  wire or_1045_nl;
  wire or_1044_nl;
  wire mux_278_nl;
  wire mux_277_nl;
  wire or_1057_nl;
  wire or_1056_nl;
  wire or_1055_nl;
  wire or_1054_nl;
  wire mux_285_nl;
  wire mux_284_nl;
  wire mux_283_nl;
  wire mux_282_nl;
  wire mux_281_nl;
  wire mux_280_nl;
  wire or_1064_nl;
  wire or_1063_nl;
  wire or_1062_nl;
  wire or_1061_nl;
  wire or_1058_nl;
  wire mux_287_nl;
  wire while_mux_1483_nl;
  wire mux_289_nl;
  wire mux_288_nl;
  wire nand_20_nl;
  wire nand_19_nl;
  wire or_1067_nl;
  wire mux_292_nl;
  wire nor_442_nl;
  wire mux_291_nl;
  wire nor_443_nl;
  wire mux_290_nl;
  wire mux_293_nl;
  wire or_1076_nl;
  wire mux_300_nl;
  wire mux_299_nl;
  wire mux_298_nl;
  wire or_1081_nl;
  wire mux_297_nl;
  wire or_1080_nl;
  wire or_1078_nl;
  wire mux_303_nl;
  wire mux_302_nl;
  wire nand_21_nl;
  wire mux_310_nl;
  wire or_1088_nl;
  wire mux_309_nl;
  wire mux_308_nl;
  wire mux_307_nl;
  wire mux_306_nl;
  wire nand_22_nl;
  wire mux_305_nl;
  wire or_1084_nl;
  wire or_1089_nl;
  wire mux_316_nl;
  wire or_1104_nl;
  wire or_1103_nl;
  wire mux_323_nl;
  wire mux_322_nl;
  wire mux_321_nl;
  wire mux_319_nl;
  wire or_1115_nl;
  wire mux_318_nl;
  wire or_1111_nl;
  wire or_1110_nl;
  wire mux_317_nl;
  wire or_1109_nl;
  wire mux_315_nl;
  wire or_1102_nl;
  wire mux_314_nl;
  wire or_1101_nl;
  wire or_1095_nl;
  wire mux_326_nl;
  wire mux_325_nl;
  wire or_1121_nl;
  wire or_1120_nl;
  wire or_1119_nl;
  wire or_1118_nl;
  wire mux_333_nl;
  wire mux_332_nl;
  wire mux_331_nl;
  wire mux_330_nl;
  wire mux_329_nl;
  wire mux_328_nl;
  wire or_1128_nl;
  wire or_1127_nl;
  wire or_1126_nl;
  wire or_1125_nl;
  wire or_1122_nl;
  wire and_580_nl;
  wire and_579_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl;
  wire weight_mem_banks_write_if_for_if_and_35_nl;
  wire weight_mem_banks_write_if_for_if_and_36_nl;
  wire weight_mem_banks_write_if_for_if_and_37_nl;
  wire weight_mem_banks_write_if_for_if_and_38_nl;
  wire weight_mem_banks_write_if_for_if_and_39_nl;
  wire weight_mem_banks_write_if_for_if_and_40_nl;
  wire weight_mem_banks_write_if_for_if_and_41_nl;
  wire weight_mem_banks_write_if_for_if_mux_7_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl;
  wire mux_123_nl;
  wire nor_461_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl;
  wire weight_mem_banks_write_if_for_if_and_28_nl;
  wire weight_mem_banks_write_if_for_if_and_29_nl;
  wire weight_mem_banks_write_if_for_if_and_30_nl;
  wire weight_mem_banks_write_if_for_if_and_31_nl;
  wire weight_mem_banks_write_if_for_if_and_32_nl;
  wire weight_mem_banks_write_if_for_if_and_33_nl;
  wire weight_mem_banks_write_if_for_if_and_34_nl;
  wire weight_mem_banks_write_if_for_if_mux_6_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl;
  wire mux_122_nl;
  wire nor_460_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl;
  wire weight_mem_banks_write_if_for_if_and_21_nl;
  wire weight_mem_banks_write_if_for_if_and_22_nl;
  wire weight_mem_banks_write_if_for_if_and_23_nl;
  wire weight_mem_banks_write_if_for_if_and_24_nl;
  wire weight_mem_banks_write_if_for_if_and_25_nl;
  wire weight_mem_banks_write_if_for_if_and_26_nl;
  wire weight_mem_banks_write_if_for_if_and_27_nl;
  wire weight_mem_banks_write_if_for_if_mux_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl;
  wire mux_121_nl;
  wire nor_459_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl;
  wire weight_mem_banks_write_if_for_if_and_14_nl;
  wire weight_mem_banks_write_if_for_if_and_15_nl;
  wire weight_mem_banks_write_if_for_if_and_16_nl;
  wire weight_mem_banks_write_if_for_if_and_17_nl;
  wire weight_mem_banks_write_if_for_if_and_18_nl;
  wire weight_mem_banks_write_if_for_if_and_19_nl;
  wire weight_mem_banks_write_if_for_if_and_20_nl;
  wire weight_mem_banks_write_if_for_if_mux_4_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl;
  wire mux_120_nl;
  wire nor_458_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl;
  wire weight_mem_banks_write_if_for_if_and_7_nl;
  wire weight_mem_banks_write_if_for_if_and_8_nl;
  wire weight_mem_banks_write_if_for_if_and_9_nl;
  wire weight_mem_banks_write_if_for_if_and_10_nl;
  wire weight_mem_banks_write_if_for_if_and_11_nl;
  wire weight_mem_banks_write_if_for_if_and_12_nl;
  wire weight_mem_banks_write_if_for_if_and_13_nl;
  wire weight_mem_banks_write_if_for_if_mux_3_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl;
  wire mux_119_nl;
  wire nor_457_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl;
  wire weight_mem_banks_write_if_for_if_and_nl;
  wire weight_mem_banks_write_if_for_if_and_1_nl;
  wire weight_mem_banks_write_if_for_if_and_2_nl;
  wire weight_mem_banks_write_if_for_if_and_3_nl;
  wire weight_mem_banks_write_if_for_if_and_4_nl;
  wire weight_mem_banks_write_if_for_if_and_5_nl;
  wire weight_mem_banks_write_if_for_if_and_6_nl;
  wire weight_mem_banks_write_if_for_if_mux_2_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl;
  wire mux_118_nl;
  wire nor_456_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_1_nl;
  wire weight_mem_banks_write_if_for_if_mux_54_nl;
  wire mux_117_nl;
  wire nor_455_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_nl;
  wire weight_mem_banks_write_if_for_if_mux_53_nl;
  wire mux_116_nl;
  wire nor_454_nl;
  wire mux1h_1_nl;
  wire[14:0] mux1h_7_nl;
  wire not_2496_nl;
  wire mux_44_nl;
  wire or_197_nl;
  wire mux_68_nl;
  wire nor_340_nl;
  wire mux_466_nl;
  wire or_1448_nl;
  wire mux_388_nl;
  wire mux_387_nl;
  wire mux_386_nl;
  wire mux_385_nl;
  wire mux_384_nl;
  wire mux_383_nl;
  wire mux_382_nl;
  wire mux_381_nl;
  wire or_1312_nl;
  wire or_1310_nl;
  wire or_1308_nl;
  wire or_1307_nl;
  wire or_1305_nl;
  wire or_1303_nl;
  wire or_1301_nl;
  wire or_1299_nl;
  wire or_1298_nl;
  wire or_1297_nl;
  wire mux_1_nl;
  wire mux_nl;
  wire nand_36_nl;
  wire nor_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [35:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_b = MUX_v_36_2_2(accum_vector_data_0_35_0_sva,
      accum_vector_data_0_35_0_sva_dfm_1_1, accum_vector_data_and_16_cse);
  wire accum_vector_data_and_17_nl;
  wire [35:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_b;
  assign accum_vector_data_and_17_nl = and_542_cse & fsm_output;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_b = MUX_v_36_2_2(accum_vector_data_7_35_0_sva,
      accum_vector_data_7_35_0_sva_dfm_1_1, accum_vector_data_and_17_nl);
  wire [35:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_b = MUX_v_36_2_2(accum_vector_data_6_35_0_sva,
      accum_vector_data_6_35_0_sva_dfm_1_1, accum_vector_data_and_16_cse);
  wire [35:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_b = MUX_v_36_2_2(accum_vector_data_5_35_0_sva,
      accum_vector_data_5_35_0_sva_dfm_1_1, accum_vector_data_and_16_cse);
  wire [35:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_b = MUX_v_36_2_2(accum_vector_data_4_35_0_sva,
      accum_vector_data_4_35_0_sva_dfm_1_1, accum_vector_data_and_16_cse);
  wire [35:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_b = MUX_v_36_2_2(accum_vector_data_3_35_0_sva,
      accum_vector_data_3_35_0_sva_dfm_1_1, accum_vector_data_and_16_cse);
  wire [35:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_b = MUX_v_36_2_2(accum_vector_data_2_35_0_sva,
      accum_vector_data_2_35_0_sva_dfm_1_1, accum_vector_data_and_16_cse);
  wire [35:0] nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_b;
  assign nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_b = MUX_v_36_2_2(accum_vector_data_1_35_0_sva,
      accum_vector_data_1_35_0_sva_dfm_1_1, accum_vector_data_and_16_cse);
  wire  nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (~ reg_rva_in_reg_rw_sva_2_cse);
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0];
  wire  nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a = PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2
      & reg_rva_in_reg_rw_sva_2_cse;
  wire [2:0] nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s = weight_write_addrs_lpi_1_dfm_1_2[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s = {(weight_read_addrs_6_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_4[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s = weight_read_addrs_7_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s = {(weight_read_addrs_2_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s = {(weight_read_addrs_4_14_2_lpi_1_dfm_1_1[0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[1:0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s = weight_read_addrs_3_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s = weight_read_addrs_5_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s = weight_read_addrs_1_lpi_1_dfm_1_1[2:0];
  wire [255:0] nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun
      = {act_port_reg_data_255_224_sva_dfm_1_1 , act_port_reg_data_223_192_sva_dfm_3
      , act_port_reg_data_191_160_sva_dfm_3 , act_port_reg_data_159_128_sva_dfm_3
      , act_port_reg_data_127_96_sva_dfm_3 , act_port_reg_data_95_64_sva_dfm_3 ,
      act_port_reg_data_63_32_sva_dfm_3 , act_port_reg_data_31_0_sva_dfm_3};
  wire [255:0] nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun
      = {rva_out_reg_data_255_240_sva_dfm_4_6 , rva_out_reg_data_239_224_sva_dfm_4_6
      , rva_out_reg_data_223_208_sva_dfm_4_6 , rva_out_reg_data_207_192_sva_dfm_4_6
      , rva_out_reg_data_191_176_sva_dfm_4_6 , rva_out_reg_data_175_160_sva_dfm_4_6
      , rva_out_reg_data_159_144_sva_dfm_4_6 , rva_out_reg_data_143_128_sva_dfm_4_6
      , rva_out_reg_data_127_112_sva_dfm_4_6 , rva_out_reg_data_111_96_sva_dfm_4_6
      , rva_out_reg_data_95_80_sva_dfm_4_6 , rva_out_reg_data_79_64_sva_dfm_4_6 ,
      rva_out_reg_data_63_sva_dfm_4_6 , rva_out_reg_data_62_48_sva_dfm_4_6 , rva_out_reg_data_47_sva_dfm_4_6
      , rva_out_reg_data_46_40_sva_dfm_4_6 , rva_out_reg_data_39_36_sva_dfm_4_6 ,
      rva_out_reg_data_35_32_sva_dfm_4_6_rsp_0 , rva_out_reg_data_35_32_sva_dfm_4_6_rsp_1
      , rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_31_mx0 , rva_out_reg_data_30_25_sva_dfm_7_5_2
      , rva_out_reg_data_30_25_sva_dfm_7_1_0 , rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_24_mx0
      , rva_out_reg_data_23_17_sva_dfm_7 , rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_16_mx0
      , rva_out_reg_data_15_9_sva_dfm_7 , rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_8_mx0
      , rva_out_reg_data_7_1_sva_dfm_7 , rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_0_mx0};
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd36),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_b[35:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd36),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_b[35:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd36),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_b[35:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd36),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_b[35:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd36),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_b[35:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd36),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_b[35:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd36),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_b[35:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_z)
    );
  PECore_mgc_mul_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd36),
  .signd_b(32'sd0),
  .width_z(32'sd43),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7 (
      .a(8'b10100111),
      .b(nl_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_b[35:0]),
      .clk(clk),
      .en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_z)
    );
  PECore_mgc_muladd1 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_cst(32'sd1),
  .signd_cst(32'sd0),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd11),
  .add_axb(32'sd1),
  .add_c(32'sd1),
  .add_d(32'sd1),
  .use_const(32'sd1)) PEManager_15U_GetWeightAddr_else_acc_4_cmp (
      .a(pe_config_output_counter_sva),
      .b(pe_manager_num_input_sva),
      .c(pe_config_input_counter_sva),
      .cst(1'b0),
      .z(PEManager_15U_GetWeightAddr_else_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_for_1_lshift_rg (
      .a(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a),
      .s(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_write_arbxbar_xbar_for_lshift_rg (
      .a(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a),
      .s(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s[2:0]),
      .z(weight_mem_write_arbxbar_xbar_for_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi PECore_PECoreRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(fsm_output)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi PECore_PECoreRun_input_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_oswt_pff(and_574_rmff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi PECore_PECoreRun_act_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(reg_act_port_Push_mioi_iswt0_cse),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun[255:0]),
      .act_port_Push_mioi_oswt_pff(and_576_cse)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi PECore_PECoreRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_oswt_pff(and_574_rmff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi PECore_PECoreRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun[255:0]),
      .rva_out_Push_mioi_oswt_pff(and_572_cse)
    );
  PECore_PECore_PECoreRun_wait_dp PECore_PECoreRun_wait_dp_inst (
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .PECoreRun_wen(PECoreRun_wen),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg(and_570_rmff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg(and_567_rmff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg(and_564_rmff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg(and_561_rmff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg(and_558_rmff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg(and_555_rmff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg(and_551_rmff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg(and_548_rmff),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo(reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_7_cse),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg(and_541_rmff),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_en),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_1(reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_1_cse),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_unreg_1(and_544_rmff),
      .PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en(PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_en),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_cgo(reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_63_cse),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg(and_535_rmff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_1(reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_40_cse),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_unreg_1(and_538_rmff)
    );
  PECore_PECore_PECoreRun_staller PECore_PECoreRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp)
    );
  PECore_PECore_PECoreRun_PECoreRun_fsm PECore_PECoreRun_PECoreRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .fsm_output(fsm_output)
    );
  assign weight_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_91);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign weight_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_91);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign weight_mem_banks_read_1_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_93);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign weight_mem_banks_read_1_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_93);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign weight_mem_banks_read_1_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_95);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 );
  assign weight_mem_banks_read_1_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_95);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign weight_mem_banks_read_1_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_97);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 );
  assign weight_mem_banks_read_1_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_97);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign weight_mem_banks_read_1_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_99);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 );
  assign weight_mem_banks_read_1_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_99);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign weight_mem_banks_read_1_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_101);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 );
  assign weight_mem_banks_read_1_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_101);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign weight_mem_banks_read_1_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_87);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 );
  assign weight_mem_banks_read_1_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_87);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign weight_mem_banks_read_1_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_89);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 );
  assign weight_mem_banks_read_1_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_89);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign weight_mem_banks_write_if_for_if_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_154);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 );
  assign weight_mem_banks_write_if_for_if_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_154);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign weight_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_155);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 );
  assign weight_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_155);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign weight_mem_banks_write_if_for_if_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_156);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 );
  assign weight_mem_banks_write_if_for_if_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_156);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1
      = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1
      = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign weight_mem_banks_read_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_157);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 );
  assign weight_mem_banks_read_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_157);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign weight_mem_banks_write_if_for_if_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_158);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 );
  assign weight_mem_banks_write_if_for_if_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_158);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2
      = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2
      = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign weight_mem_banks_read_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_159);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 );
  assign weight_mem_banks_read_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_159);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign weight_mem_banks_write_if_for_if_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_160);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 );
  assign weight_mem_banks_write_if_for_if_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_160);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3
      = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3
      = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign weight_mem_banks_read_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_161);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 );
  assign weight_mem_banks_read_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_161);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign weight_mem_banks_write_if_for_if_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_162);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 );
  assign weight_mem_banks_write_if_for_if_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_162);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4
      = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4
      = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign weight_mem_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_163);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 );
  assign weight_mem_banks_read_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_163);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign weight_mem_banks_write_if_for_if_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_164);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 );
  assign weight_mem_banks_write_if_for_if_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_164);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5
      = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5
      = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign weight_mem_banks_read_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_165);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 );
  assign weight_mem_banks_read_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_165);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign weight_mem_banks_write_if_for_if_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_166);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 );
  assign weight_mem_banks_write_if_for_if_mux_33_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_166);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6
      = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6
      = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign weight_mem_banks_read_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_167);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 );
  assign weight_mem_banks_read_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_167);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign weight_mem_banks_write_if_for_if_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_168);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 );
  assign weight_mem_banks_write_if_for_if_mux_37_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_168);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7
      = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7
      = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign weight_mem_banks_read_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_169);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 );
  assign weight_mem_banks_read_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_169);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign input_mem_banks_write_1_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_179);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 );
  assign input_mem_banks_write_1_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_179);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8
      = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_3 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8
      = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign input_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_176);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 );
  assign input_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_176);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign input_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_188);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 );
  assign input_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_188);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9
      = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_1 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9
      = input_mem_banks_write_if_for_if_mux_1_cse;
  assign input_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_191);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 );
  assign input_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_191);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign and_535_rmff = (((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_8 & while_stage_0_10) | and_dcpl_532
      | and_dcpl_530) & fsm_output;
  assign and_538_rmff = (and_537_cse | and_dcpl_532 | and_dcpl_530) & fsm_output;
  assign and_540_nl = or_tmp_75 & or_tmp_76;
  assign nor_18_nl = ~(PECore_RunMac_PECore_RunMac_if_and_svs_st_10 | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_10));
  assign mux_70_nl = MUX_s_1_2_2(or_tmp_75, and_540_nl, nor_18_nl);
  assign and_541_rmff = (~ mux_70_nl) & fsm_output;
  assign or_697_nl = (~ while_stage_0_10) | PECore_RunMac_PECore_RunMac_if_and_svs_st_8
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  assign and_543_nl = or_tmp_78 & (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 |
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign mux_71_nl = MUX_s_1_2_2(or_tmp_78, and_543_nl, while_stage_0_10);
  assign and_988_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9 & while_stage_0_11;
  assign mux_72_nl = MUX_s_1_2_2(or_697_nl, mux_71_nl, and_988_nl);
  assign mux_73_nl = MUX_s_1_2_2(or_tmp_75, mux_72_nl, PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8);
  assign and_544_rmff = (~ mux_73_nl) & fsm_output;
  assign or_700_nl = (while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_336_itm_1) & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3)
      | and_tmp_2;
  assign nand_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~((~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_336_itm_1 | (~
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3)))
      | and_tmp_2)));
  assign mux_75_nl = MUX_s_1_2_2(and_tmp_2, nand_nl, while_stage_0_7);
  assign mux_76_nl = MUX_s_1_2_2(or_700_nl, mux_75_nl, weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign and_548_rmff = (mux_76_nl | and_dcpl_544) & fsm_output;
  assign or_706_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | and_tmp_3;
  assign or_705_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3;
  assign or_704_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_1 | weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3;
  assign mux_78_nl = MUX_s_1_2_2(or_705_nl, or_704_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_79_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3,
      mux_78_nl, while_stage_0_6);
  assign mux_80_nl = MUX_s_1_2_2(or_706_nl, mux_79_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_81_nl = MUX_s_1_2_2(and_tmp_3, mux_80_nl, while_stage_0_7);
  assign or_703_nl = (~((~ while_stage_0_7) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)))
      | and_tmp_3;
  assign mux_82_nl = MUX_s_1_2_2(mux_81_nl, or_703_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_328_itm_1);
  assign and_551_rmff = (mux_82_nl | and_dcpl_546) & fsm_output;
  assign or_710_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_4;
  assign or_709_nl = (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2)))
      | and_tmp_4;
  assign mux_84_nl = MUX_s_1_2_2(or_710_nl, or_709_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_85_nl = MUX_s_1_2_2(and_tmp_4, mux_84_nl, while_stage_0_6);
  assign and_555_rmff = (mux_85_nl | and_dcpl_164) & fsm_output;
  assign or_718_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_5;
  assign or_1149_nl = (~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_1)) | and_tmp_5;
  assign mux_87_nl = MUX_s_1_2_2(or_718_nl, or_1149_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_88_nl = MUX_s_1_2_2(and_tmp_5, mux_87_nl, while_stage_0_6);
  assign and_558_rmff = (mux_88_nl | and_dcpl_162) & fsm_output;
  assign or_722_nl = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_6;
  assign or_1150_nl = (~((~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1)) | and_tmp_6;
  assign mux_90_nl = MUX_s_1_2_2(or_722_nl, or_1150_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_91_nl = MUX_s_1_2_2(and_tmp_6, mux_90_nl, while_stage_0_6);
  assign and_561_rmff = (mux_91_nl | and_dcpl_160) & fsm_output;
  assign or_726_nl = (while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1) & reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse)
      | and_tmp_7;
  assign nand_3_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (~((~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1 | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse)))
      | and_tmp_7)));
  assign mux_93_nl = MUX_s_1_2_2(and_tmp_7, nand_3_nl, while_stage_0_6);
  assign mux_94_nl = MUX_s_1_2_2(or_726_nl, mux_93_nl, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign and_564_rmff = (mux_94_nl | and_dcpl_158) & fsm_output;
  assign or_735_nl = (while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1) & reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse)
      | and_tmp_8;
  assign nand_4_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (~((~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1 | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse)))
      | and_tmp_8)));
  assign mux_97_nl = MUX_s_1_2_2(and_tmp_8, nand_4_nl, while_stage_0_6);
  assign mux_98_nl = MUX_s_1_2_2(or_735_nl, mux_97_nl, weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign and_567_rmff = (mux_98_nl | and_dcpl_156) & fsm_output;
  assign or_739_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | and_tmp_9;
  assign or_1151_nl = (~((~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1)) | and_tmp_9;
  assign mux_100_nl = MUX_s_1_2_2(or_739_nl, or_1151_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_101_nl = MUX_s_1_2_2(and_tmp_9, mux_100_nl, while_stage_0_6);
  assign and_570_rmff = (mux_101_nl | and_dcpl_154) & fsm_output;
  assign and_1065_itm = PECore_UpdateFSM_switch_lp_nor_7_itm_1 & PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      & pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign and_756_itm = pe_config_is_zero_first_sva & PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      & pe_manager_zero_active_sva;
  assign and_768_cse = PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign mux_467_nl = MUX_s_1_2_2(and_1065_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_756_itm);
  assign and_767_nl = start_PopNB_mioi_data_rsc_z_mxwt & start_PopNB_mioi_return_rsc_z_mxwt
      & PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign mux_110_nl = MUX_s_1_2_2(mux_467_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_767_nl);
  assign mux_349_nl = MUX_s_1_2_2(and_1065_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_756_itm);
  assign mux_106_nl = MUX_s_1_2_2(mux_349_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_768_cse);
  assign mux_111_nl = MUX_s_1_2_2(mux_110_nl, mux_106_nl, or_142_cse);
  assign mux_469_nl = MUX_s_1_2_2(and_1065_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_756_itm);
  assign mux_468_nl = MUX_s_1_2_2(mux_469_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_768_cse);
  assign or_140_nl = pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]);
  assign mux_107_nl = MUX_s_1_2_2(mux_468_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_140_nl);
  assign or_139_nl = (state_2_1_sva!=2'b10) | state_0_sva;
  assign mux_108_nl = MUX_s_1_2_2(mux_107_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_139_nl);
  assign mux_109_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_nor_7_itm_1, mux_108_nl,
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign mux_112_nl = MUX_s_1_2_2(mux_111_nl, mux_109_nl, PECore_UpdateFSM_switch_lp_equal_tmp_5_1);
  assign mux_113_nl = MUX_s_1_2_2(mux_112_nl, state_0_sva, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_114_nl = MUX_s_1_2_2(or_142_cse, mux_113_nl, while_stage_0_3);
  assign or_138_nl = while_stage_0_3 | (state_2_1_sva!=2'b00) | state_0_sva;
  assign or_137_nl = (state_2_1_sva_dfm_1!=2'b00);
  assign mux_115_cse = MUX_s_1_2_2(mux_114_nl, or_138_nl, or_137_nl);
  assign and_574_rmff = (~ mux_115_cse) & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign PECore_DecodeAxiRead_switch_lp_and_2_cse = PECoreRun_wen & and_dcpl_8;
  assign rva_out_reg_data_and_26_cse = PECoreRun_wen & and_dcpl_8 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_10) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10)
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 | rva_in_reg_rw_sva_st_10));
  assign rva_out_reg_data_and_191_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_15_9_sva_dfm_10_enexo;
  assign rva_out_reg_data_and_192_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_23_17_sva_dfm_8_enexo;
  assign rva_out_reg_data_and_29_cse = PECoreRun_wen & and_dcpl_7;
  assign rva_out_reg_data_and_193_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_255_240_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_194_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_239_224_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_195_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_223_208_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_196_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_207_192_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_197_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_191_176_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_198_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_175_160_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_199_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_159_144_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_200_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_143_128_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_201_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_127_112_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_202_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_111_96_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_203_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_95_80_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_204_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_205_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_79_64_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_206_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_5_enexo;
  assign rva_out_reg_data_and_207_enex5 = rva_out_reg_data_and_29_cse & reg_rva_out_reg_data_62_48_sva_dfm_4_5_enexo;
  assign input_mem_banks_read_read_data_and_cse = PECoreRun_wen & and_dcpl_7 & (~
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8) & input_read_req_valid_lpi_1_dfm_1_10;
  assign weight_port_read_out_data_and_125_cse = PECoreRun_wen & and_dcpl_6 & (~
      rva_in_reg_rw_sva_st_1_10) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8;
  assign weight_port_read_out_data_and_172_enex5 = weight_port_read_out_data_and_125_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_cse = PECoreRun_wen & (~((~(while_stage_0_13 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11))
      | rva_in_reg_rw_sva_11));
  assign input_mem_banks_read_read_data_and_57_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5_enexo;
  assign input_mem_banks_read_read_data_and_58_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5_enexo;
  assign weight_port_read_out_data_and_173_enex5 = weight_port_read_out_data_and_125_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_5_1_enexo;
  assign input_mem_banks_read_read_data_and_59_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5_enexo;
  assign input_mem_banks_read_read_data_and_60_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5_enexo;
  assign rva_in_reg_rw_and_cse = PECoreRun_wen & while_stage_0_12;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_cse = PECoreRun_wen & and_dcpl_6
      & (~(rva_in_reg_rw_sva_st_1_10 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8))
      & (~(rva_in_reg_rw_sva_10 | input_read_req_valid_lpi_1_dfm_1_10)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9;
  assign PECore_PushOutput_if_and_cse = PECoreRun_wen & and_dcpl_24;
  assign and_1072_cse = ((PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11))
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_11) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11)
      & while_stage_0_13 & PECoreRun_wen;
  assign accum_vector_data_and_cse = PECoreRun_wen & (~ or_tmp_76);
  assign accum_vector_data_and_24_enex5 = accum_vector_data_and_cse & reg_accum_vector_data_6_35_0_sva_dfm_1_1_enexo;
  assign accum_vector_data_and_25_enex5 = accum_vector_data_and_cse & reg_accum_vector_data_5_35_0_sva_dfm_1_1_enexo;
  assign accum_vector_data_and_26_enex5 = accum_vector_data_and_cse & reg_accum_vector_data_4_35_0_sva_dfm_1_1_enexo;
  assign accum_vector_data_and_27_enex5 = accum_vector_data_and_cse & reg_accum_vector_data_3_35_0_sva_dfm_1_1_enexo;
  assign accum_vector_data_and_28_enex5 = accum_vector_data_and_cse & reg_accum_vector_data_2_35_0_sva_dfm_1_1_enexo;
  assign accum_vector_data_and_29_enex5 = accum_vector_data_and_cse & reg_accum_vector_data_1_35_0_sva_dfm_1_1_enexo;
  assign accum_vector_data_and_30_enex5 = accum_vector_data_and_cse & reg_accum_vector_data_0_35_0_sva_dfm_1_1_enexo;
  assign PECore_RunMac_if_and_1_cse = PECoreRun_wen & and_542_cse;
  assign and_1099_cse = ((~ while_stage_0_12) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_10
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_9 | PECore_UpdateFSM_switch_lp_equal_tmp_2_9)
      & while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9)
      & PECoreRun_wen;
  assign while_if_and_6_cse = PECoreRun_wen & while_stage_0_11;
  assign accum_vector_data_and_7_enex5 = PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9
      | (~ while_stage_0_11))) & reg_accum_vector_data_7_35_0_sva_dfm_1_1_enexo;
  assign PECore_RunMac_if_and_2_cse = PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & while_stage_0_10;
  assign while_if_and_7_cse = PECoreRun_wen & while_stage_0_10;
  assign PECore_RunMac_if_and_3_cse = PECoreRun_wen & (and_dcpl_40 | and_dcpl_344);
  assign while_if_and_8_cse = PECoreRun_wen & while_stage_0_9;
  assign PECore_RunMac_if_and_4_cse = PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & rva_in_reg_rw_sva_st_1_6)) & while_stage_0_8;
  assign while_if_and_9_cse = PECoreRun_wen & while_stage_0_8;
  assign input_mem_banks_read_1_read_data_and_cse = PECoreRun_wen & and_537_cse;
  assign input_mem_banks_read_1_read_data_and_5_enex5 = input_mem_banks_read_1_read_data_and_cse
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  assign weight_mem_run_3_for_5_and_163_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_162_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign or_1189_cse = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~ while_stage_0_8);
  assign weight_port_read_out_data_and_enex5 = PECoreRun_wen & (~(or_1189_cse | (~
      weight_mem_run_3_for_land_2_lpi_1_dfm_3))) & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000;
  assign weight_mem_run_3_for_aelse_and_cse = PECoreRun_wen & while_stage_0_7;
  assign weight_port_read_out_data_and_1_cse = PECoreRun_wen & (~(or_1189_cse | (~
      weight_mem_run_3_for_land_3_lpi_1_dfm_3)));
  assign weight_port_read_out_data_and_174_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000;
  assign data_in_tmp_operator_2_for_and_1_cse = PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & weight_mem_run_3_for_land_3_lpi_1_dfm_2 & while_stage_0_7;
  assign weight_port_read_out_data_and_175_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000001;
  assign weight_port_read_out_data_and_176_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000002;
  assign weight_port_read_out_data_and_177_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000003;
  assign weight_port_read_out_data_and_178_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000004;
  assign weight_port_read_out_data_and_179_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000005;
  assign weight_port_read_out_data_and_180_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000006;
  assign weight_port_read_out_data_and_181_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000007;
  assign weight_port_read_out_data_and_182_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000008;
  assign weight_port_read_out_data_and_183_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000009;
  assign weight_port_read_out_data_and_184_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000010;
  assign weight_port_read_out_data_and_185_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000011;
  assign weight_port_read_out_data_and_186_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000012;
  assign weight_port_read_out_data_and_187_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000013;
  assign weight_port_read_out_data_and_188_enex5 = weight_port_read_out_data_and_1_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000014;
  assign weight_port_read_out_data_and_16_cse = PECoreRun_wen & (~(or_1189_cse |
      (~ weight_mem_run_3_for_land_5_lpi_1_dfm_3)));
  assign weight_port_read_out_data_and_189_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000;
  assign data_in_tmp_operator_2_for_and_16_cse = PECoreRun_wen & and_dcpl_45 & weight_mem_run_3_for_land_5_lpi_1_dfm_2;
  assign weight_port_read_out_data_and_190_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000001;
  assign weight_port_read_out_data_and_191_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000002;
  assign weight_port_read_out_data_and_192_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000003;
  assign weight_port_read_out_data_and_193_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000004;
  assign weight_port_read_out_data_and_194_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000005;
  assign weight_port_read_out_data_and_195_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000006;
  assign weight_port_read_out_data_and_196_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000007;
  assign weight_port_read_out_data_and_197_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000008;
  assign weight_port_read_out_data_and_198_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000009;
  assign weight_port_read_out_data_and_199_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000010;
  assign weight_port_read_out_data_and_200_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000011;
  assign weight_port_read_out_data_and_201_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000012;
  assign weight_port_read_out_data_and_202_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000013;
  assign weight_port_read_out_data_and_203_enex5 = weight_port_read_out_data_and_16_cse
      & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000014;
  assign weight_port_read_out_data_and_31_enex5 = PECoreRun_wen & (~(or_1189_cse
      | (~ weight_mem_run_3_for_land_4_lpi_1_dfm_3))) & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000;
  assign PECore_RunMac_if_and_5_cse = PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & rva_in_reg_rw_sva_st_1_5)) & while_stage_0_7;
  assign rva_in_reg_rw_and_2_cse = PECoreRun_wen & and_dcpl_56;
  assign input_mem_banks_read_1_read_data_and_1_enex5 = PECoreRun_wen & and_dcpl_57
      & reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  assign PECore_RunMac_if_and_6_cse = PECoreRun_wen & and_dcpl_57;
  assign weight_port_read_out_data_7_15_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[255:240]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[255:240]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[239:224]), weight_port_read_out_data_7_15_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_143_itm_1 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign nor_500_cse = ~((weight_read_addrs_7_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_356_nl = MUX_s_1_2_2((weight_read_addrs_7_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_7_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_7_lpi_1_dfm_3_2_0[0]);
  assign mux_357_nl = MUX_s_1_2_2(mux_356_nl, nor_500_cse, weight_read_addrs_7_lpi_1_dfm_3_2_0[2]);
  assign and_1130_cse = (mux_357_nl | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_port_read_out_data_7_14_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[239:224]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[239:224]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[223:208]), weight_port_read_out_data_7_14_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_132_itm_1 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_asn_451 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign xor_1_cse = (weight_read_addrs_7_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[2]);
  assign and_1135_cse = (xor_1_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_port_read_out_data_7_13_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[223:208]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[223:208]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[207:192]), weight_port_read_out_data_7_13_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_asn_451 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign and_1141_cse = (and_1135_cse | or_dcpl_761 | weight_mem_run_3_for_5_and_140_itm_2)
      & and_dcpl_808 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign weight_port_read_out_data_7_12_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[207:192]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[207:192]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[191:176]), weight_port_read_out_data_7_12_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_132_itm_1 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_11_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[191:176]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[191:176]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[175:160]), weight_port_read_out_data_7_11_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_asn_451 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_10_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[175:160]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[175:160]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[159:144]), weight_port_read_out_data_7_10_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_143_itm_1 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign and_1156_cse = (and_1130_cse | or_dcpl_753 | or_dcpl_774) & and_dcpl_808
      & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign weight_port_read_out_data_7_9_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[159:144]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[159:144]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[143:128]), weight_port_read_out_data_7_9_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_143_itm_1 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_8_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[143:128]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[143:128]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[127:112]), weight_port_read_out_data_7_8_sva_dfm_1,
      {weight_mem_run_3_for_5_and_153 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_143_itm_1 , weight_mem_run_3_for_5_asn_451 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign and_1165_cse = (xor_1_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_port_read_out_data_7_7_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[111:96]), weight_port_read_out_data_7_7_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_asn_451 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_6_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[95:80]), weight_port_read_out_data_7_6_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_143_itm_1 , weight_mem_run_3_for_5_asn_451 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_5_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[79:64]), weight_port_read_out_data_7_5_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_142_itm_1
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_4_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[63:48]), weight_port_read_out_data_7_4_sva_dfm_1,
      {weight_mem_run_3_for_5_and_153 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_132_itm_1 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_143_itm_1 , weight_mem_run_3_for_5_asn_451 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_3_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[47:32]), weight_port_read_out_data_7_3_sva_dfm_1,
      {weight_mem_run_3_for_5_and_153 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_132_itm_1 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_asn_451 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_2_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[31:16]), weight_port_read_out_data_7_2_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_132_itm_1 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_1_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[15:0]), weight_port_read_out_data_7_1_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign and_1201_cse = (and_1130_cse | or_dcpl_766 | or_dcpl_774) & and_dcpl_808
      & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign weight_port_read_out_data_7_0_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]),
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9, weight_port_read_out_data_7_0_sva_dfm_1,
      {weight_mem_run_3_for_5_and_157 , weight_mem_run_3_for_5_asn_445 , weight_mem_run_3_for_5_asn_447
      , weight_mem_run_3_for_5_and_140_itm_2 , weight_mem_run_3_for_5_asn_449 , weight_mem_run_3_for_5_and_126_itm_2
      , weight_mem_run_3_for_5_and_135_itm_2 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_mem_run_3_for_aelse_and_5_cse = PECoreRun_wen & while_stage_0_6;
  assign weight_port_read_out_data_5_15_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[255:240]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[255:240]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[239:224]), weight_port_read_out_data_5_15_sva_dfm_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_453
      , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_1_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign nor_508_cse = ~((weight_read_addrs_5_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_372_nl = MUX_s_1_2_2((weight_read_addrs_5_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_5_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_5_lpi_1_dfm_3_2_0[0]);
  assign mux_373_nl = MUX_s_1_2_2(mux_372_nl, nor_508_cse, weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign and_1210_cse = (mux_373_nl | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_port_read_out_data_5_14_sva_dfm_3 = MUX1HOT_v_16_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[239:224]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[239:224]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[223:208]), weight_port_read_out_data_5_14_sva_dfm_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_453
      , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_6_itm_1_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign or_1284_cse = (~ while_stage_0_6) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign weight_read_addrs_and_2_enex5 = PECoreRun_wen & ((weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
      & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]))) | (weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
      & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6])))) & and_dcpl_76 &
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse = PECoreRun_wen & and_dcpl_87;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse
      & (reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo);
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse = PECoreRun_wen & and_dcpl_89;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse
      & (reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo_1
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3_enexo
      | reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo_1);
  assign while_if_and_12_cse = PECoreRun_wen & while_stage_0_5;
  assign weight_mem_read_arbxbar_arbiters_next_and_cse = PECoreRun_wen & fsm_output;
  assign weight_mem_read_arbxbar_arbiters_next_and_52_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((nor_276_cse & (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) |
      (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]))) & nor_279_cse) | or_188_cse);
  assign weight_mem_read_arbxbar_arbiters_next_and_58_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_115_cse | or_188_cse);
  assign weight_mem_read_arbxbar_arbiters_next_and_64_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & or_dcpl_47;
  assign weight_mem_read_arbxbar_arbiters_next_and_69_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & or_dcpl_48;
  assign weight_mem_read_arbxbar_arbiters_next_and_74_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & or_dcpl_50;
  assign weight_mem_read_arbxbar_arbiters_next_and_79_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (or_188_cse | (~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp));
  assign weight_mem_read_arbxbar_arbiters_next_and_85_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & or_dcpl_53;
  assign weight_mem_read_arbxbar_arbiters_next_and_90_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4));
  assign weight_read_addrs_and_4_cse = PECoreRun_wen & (and_dcpl_130 | and_dcpl_129
      | and_dcpl_128 | and_dcpl_127 | and_dcpl_126 | and_dcpl_125 | and_dcpl_124
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | and_dcpl_123) & while_stage_0_4;
  assign weight_write_data_data_and_cse = PECoreRun_wen & and_dcpl_133 & ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7:6]!=2'b00));
  assign weight_write_data_data_and_48_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_49_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_50_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_51_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_52_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_53_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_54_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_55_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_56_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_57_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_58_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_59_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_60_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_61_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_62_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_63_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_addrs_and_enex5 = weight_write_data_data_and_cse & reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  assign weight_mem_write_arbxbar_xbar_for_1_for_and_cse = PECoreRun_wen & and_dcpl_133;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
      = PECoreRun_wen & and_dcpl_137;
  assign PECore_RunFSM_switch_lp_and_cse = PECoreRun_wen & while_stage_0_4;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_5_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 & and_dcpl_137;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse
      = PECoreRun_wen & and_dcpl_137 & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse
      = PECoreRun_wen & or_185_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign Arbiter_8U_Roundrobin_pick_1_and_15_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8
      & and_dcpl_137;
  assign Arbiter_8U_Roundrobin_pick_and_85_cse = PECoreRun_wen & (while_stage_0_4
      | and_dcpl_590) & fsm_output & or_188_cse;
  assign Arbiter_8U_Roundrobin_pick_1_and_22_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9
      & and_dcpl_137;
  assign Arbiter_8U_Roundrobin_pick_1_and_64_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign weight_write_data_data_and_16_cse = PECoreRun_wen & and_dcpl_172;
  assign weight_write_data_data_and_64_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_65_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_66_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_67_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_68_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_69_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_70_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_71_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_72_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_73_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_74_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_75_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_76_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_77_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_78_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_79_enex5 = weight_write_data_data_and_16_cse
      & reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  assign weight_write_addrs_and_3_enex5 = weight_write_data_data_and_16_cse & reg_weight_write_addrs_lpi_1_dfm_1_1_enexo;
  assign rva_in_reg_rw_and_3_cse = PECoreRun_wen & while_stage_0_3;
  assign weight_read_addrs_and_enex5 = weight_write_data_data_and_16_cse & reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  assign state_and_cse = weight_mem_read_arbxbar_arbiters_next_and_cse & nand_83_cse;
  assign nor_521_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:14]!=2'b00));
  assign nor_518_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10:8]!=3'b000));
  assign nor_520_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:11]!=3'b000));
  assign and_1227_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & while_stage_0_3;
  assign pe_config_num_manager_and_cse = PECoreRun_wen & (~(or_dcpl_649 | or_dcpl_648
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~(PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])))));
  assign rva_in_reg_rw_and_4_cse = PECoreRun_wen & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign PECore_UpdateFSM_switch_lp_and_9_cse = PECoreRun_wen & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign or_142_cse = (state_2_1_sva!=2'b00) | state_0_sva;
  assign or_1293_cse = (~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]!=2'b00) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]!=2'b01);
  assign nor_523_cse = ~((~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1);
  assign and_1437_cse = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  assign pe_config_UpdateManagerCounter_if_if_and_enex5 = PECoreRun_wen & reg_pe_config_num_output_enexo;
  assign PECore_DecodeAxiRead_switch_lp_and_cse = PECoreRun_wen & (~(nand_83_cse
      | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
  assign PECore_DecodeAxiWrite_switch_lp_and_cse = PECoreRun_wen & (~ or_dcpl_648);
  assign PECore_UpdateFSM_switch_lp_and_16_cse = PECoreRun_wen & and_dcpl_40;
  assign weight_port_read_out_data_and_131_cse = PECoreRun_wen & and_dcpl_195;
  assign nand_72_cse = ~(while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6);
  assign nor_526_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]) | (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]));
  assign mux_391_nl = MUX_s_1_2_2((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]),
      (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])), reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign mux_392_nl = MUX_s_1_2_2(mux_391_nl, nor_526_cse, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]);
  assign or_1318_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1
      | mux_392_nl;
  assign mux_393_nl = MUX_s_1_2_2(nand_72_cse, or_1318_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_1266_cse = (mux_393_nl | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1) & and_dcpl_195
      & PECoreRun_wen;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2:1]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1:0]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_or_3_cse = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) & nor_526_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]) & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_1017_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_28 & (~ or_dcpl);
  assign and_1018_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_3_cse & (~
      or_dcpl);
  assign and_1019_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      & (~ or_dcpl);
  assign and_1020_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1
      & (~ or_dcpl);
  assign and_1021_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_itm_1
      & (~ or_dcpl);
  assign and_1022_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1
      & (~ or_dcpl);
  assign nor_472_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl);
  assign weight_read_addrs_and_15_cse = PECoreRun_wen & while_stage_0_6 & weight_mem_run_3_for_land_5_lpi_1_dfm_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_read_addrs_and_16_cse = PECoreRun_wen & weight_mem_run_3_for_land_7_lpi_1_dfm_1
      & while_stage_0_6 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_port_read_out_data_and_50_cse = PECoreRun_wen & (while_and_1256_cse
      | while_and_46_tmp) & while_stage_0_7;
  assign weight_port_read_out_data_and_134_cse = PECoreRun_wen & weight_mem_run_3_for_land_7_lpi_1_dfm_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7 & fsm_output & ((~(weight_mem_run_3_for_land_7_lpi_1_dfm_1
      & while_stage_0_6)) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_port_read_out_data_and_78_cse = PECoreRun_wen & (~(or_dcpl_633 |
      (~ weight_mem_run_3_for_land_2_lpi_1_dfm_2)));
  assign nor_273_nl = ~((~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp));
  assign mux_2_nl = MUX_s_1_2_2(nor_273_nl, weight_mem_run_3_for_land_6_lpi_1_dfm_1,
      while_stage_0_6);
  assign or_8_nl = while_stage_0_6 | (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp);
  assign mux_3_nl = MUX_s_1_2_2((~ mux_2_nl), or_8_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_port_read_out_data_and_150_cse = PECoreRun_wen & (~(or_dcpl_633 |
      (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2) | (~ fsm_output))) & mux_3_nl;
  assign weight_port_read_out_data_and_109_cse = PECoreRun_wen & (~(or_dcpl_633 |
      (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)));
  assign and_1441_cse = weight_mem_run_3_for_land_1_lpi_1_dfm_3 & weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_6_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_374_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1 & while_stage_0_6 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_378_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1 & while_stage_0_6 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_382_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_4_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_387_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1 & while_stage_0_6 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_389_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_2_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse = PECoreRun_wen & while_stage_0_6
      & weight_mem_run_3_for_land_1_lpi_1_dfm_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_read_addrs_and_19_cse = PECoreRun_wen & and_dcpl_85;
  assign or_188_cse = (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign or_185_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
      = weight_mem_read_arbxbar_arbiters_next_and_cse & or_188_cse;
  assign weight_read_addrs_and_27_enex5 = weight_write_data_data_and_16_cse & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  assign operator_15_false_1_and_cse = PECoreRun_wen & (~(and_dcpl_588 | or_188_cse));
  assign PEManager_15U_PEManagerWrite_and_enex5 = PECoreRun_wen & reg_rva_in_reg_rw_sva_st_1_1_cse
      & (~ PECore_DecodeAxiWrite_switch_lp_equal_tmp_2) & (~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1)) & PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_in_reg_data_sva_1_enexo;
  assign pe_manager_num_input_and_cse = PECoreRun_wen & (~(or_dcpl_649 | nand_83_cse
      | or_dcpl_700));
  assign pe_config_is_valid_and_cse = PECoreRun_wen & (~(PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1
      | PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (~ nand_83_cse);
  assign nor_534_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:6]!=2'b00));
  assign and_1294_cse = (((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5:2]==4'b0000)
      & nor_534_cse & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:8]==6'b000000) &
      nor_521_cse & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]==2'b01)) | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | (~(reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3))) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01)
      & rva_in_PopNB_mioi_return_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]==2'b00)
      & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & rva_in_reg_rw_and_4_cse;
  assign while_if_and_16_cse = PECoreRun_wen & and_dcpl_180;
  assign rva_in_reg_rw_and_5_cse = PECoreRun_wen & and_dcpl_76;
  assign rva_in_reg_rw_and_6_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9
      & while_stage_0_11;
  assign input_mem_banks_read_read_data_and_9_cse = PECoreRun_wen & and_dcpl_231
      & input_read_req_valid_lpi_1_dfm_1_9 & while_stage_0_11;
  assign input_mem_banks_read_read_data_and_61_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo;
  assign input_mem_banks_read_read_data_and_62_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo;
  assign input_mem_banks_read_read_data_and_63_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo;
  assign input_mem_banks_read_read_data_and_64_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse = PECoreRun_wen & and_dcpl_230
      & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 | input_read_req_valid_lpi_1_dfm_1_9))
      & (~ rva_in_reg_rw_sva_9) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 &
      while_stage_0_11;
  assign input_mem_banks_read_1_read_data_and_2_enex5 = PECoreRun_wen & PECore_RunMac_PECore_RunMac_if_and_svs_st_3
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  assign input_read_req_valid_and_1_cse = PECoreRun_wen & and_dcpl_230 & while_stage_0_11;
  assign PECore_DecodeAxiRead_switch_lp_and_7_cse = PECoreRun_wen & and_dcpl_231
      & and_dcpl_241 & while_stage_0_11;
  assign rva_out_reg_data_and_47_cse = PECoreRun_wen & and_dcpl_231 & and_dcpl_241
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_9) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8
      & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9)
      & (~ rva_in_reg_rw_sva_st_9) & while_stage_0_11;
  assign rva_out_reg_data_and_208_enex5 = rva_out_reg_data_and_47_cse & reg_rva_out_reg_data_30_25_sva_dfm_7_enexo;
  assign rva_out_reg_data_and_209_enex5 = rva_out_reg_data_and_47_cse & reg_rva_out_reg_data_23_17_sva_dfm_7_enexo;
  assign rva_out_reg_data_and_210_enex5 = rva_out_reg_data_and_47_cse & reg_rva_out_reg_data_15_9_sva_dfm_9_enexo;
  assign weight_port_read_out_data_and_164_cse = PECoreRun_wen & and_dcpl_230 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7
      & while_stage_0_11;
  assign weight_port_read_out_data_and_204_enex5 = weight_port_read_out_data_and_164_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_4_enexo;
  assign rva_out_reg_data_and_211_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_212_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_213_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_62_48_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_214_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_255_240_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_215_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_239_224_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_216_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_223_208_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_217_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_207_192_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_218_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_191_176_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_219_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_175_160_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_220_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_159_144_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_221_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_143_128_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_222_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_127_112_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_223_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_111_96_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_224_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_95_80_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_225_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_79_64_sva_dfm_4_4_enexo;
  assign weight_mem_banks_load_store_for_else_and_cse = PECoreRun_wen & and_dcpl_253
      & and_dcpl_56;
  assign weight_mem_banks_load_store_for_else_and_72_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1 & and_dcpl_56;
  assign and_1025_cse = nor_335_cse & (~ or_dcpl_719);
  assign and_1026_cse = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])
      & (~ or_dcpl_719);
  assign and_1027_cse = and_dcpl_657 & (~ or_dcpl_719);
  assign mux_42_nl = MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]),
      (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign nor_291_nl = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]!=2'b00));
  assign mux_43_nl = MUX_s_1_2_2(mux_42_nl, nor_291_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign weight_mem_banks_load_store_for_else_and_73_cse = PECoreRun_wen & mux_43_nl
      & and_dcpl_258 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign weight_mem_banks_load_store_for_else_and_74_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1
      & while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign weight_mem_banks_load_store_for_else_and_75_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1
      & while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_248_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[31:16]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_248_nl);
  assign nor_335_cse = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2:1]!=2'b00));
  assign weight_read_addrs_and_23_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse
      & and_dcpl_274;
  assign and_279_cse = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) & PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp;
  assign rva_in_reg_rw_and_9_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
      & while_stage_0_10;
  assign pe_manager_base_weight_and_5_cse = PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_7_or_cse
      & and_dcpl_274;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_396_cse = PECoreRun_wen
      & (weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_398_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_402_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_159_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_163_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_1_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign input_mem_banks_read_read_data_and_18_cse = PECoreRun_wen & and_dcpl_313
      & input_read_req_valid_lpi_1_dfm_1_8 & while_stage_0_10;
  assign input_mem_banks_read_read_data_and_65_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_66_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_67_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo;
  assign input_mem_banks_read_read_data_and_68_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse = PECoreRun_wen & and_dcpl_312
      & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 | rva_in_reg_rw_sva_8))
      & (~ input_read_req_valid_lpi_1_dfm_1_8) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7
      & while_stage_0_10;
  assign PECore_UpdateFSM_switch_lp_and_18_cse = PECoreRun_wen & and_dcpl_320;
  assign input_mem_banks_read_1_read_data_and_3_enex5 = PECoreRun_wen & and_dcpl_321
      & while_stage_0_4 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  assign input_read_req_valid_and_2_cse = PECoreRun_wen & and_dcpl_312 & while_stage_0_10;
  assign PECore_DecodeAxiRead_switch_lp_and_11_cse = PECoreRun_wen & and_dcpl_313
      & and_dcpl_325 & while_stage_0_10;
  assign rva_out_reg_data_and_68_cse = PECoreRun_wen & and_dcpl_313 & and_dcpl_325
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_8) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7
      & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8)
      & while_stage_0_10 & (~ rva_in_reg_rw_sva_st_8);
  assign rva_out_reg_data_and_226_enex5 = rva_out_reg_data_and_68_cse & reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_227_enex5 = rva_out_reg_data_and_68_cse & reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  assign weight_port_read_out_data_and_166_cse = PECoreRun_wen & and_dcpl_312 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6
      & while_stage_0_10;
  assign weight_port_read_out_data_and_205_enex5 = weight_port_read_out_data_and_166_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_228_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_229_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_230_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_62_48_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_231_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_255_240_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_232_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_239_224_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_233_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_223_208_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_234_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_207_192_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_235_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_191_176_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_236_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_175_160_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_237_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_159_144_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_238_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_143_128_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_239_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_127_112_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_240_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_111_96_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_241_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_95_80_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_242_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_79_64_sva_dfm_4_3_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_7_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_125_tmp;
  assign weight_mem_write_arbxbar_xbar_for_empty_and_3_enex5 = rva_in_reg_rw_and_5_cse
      & reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  assign PECore_RunMac_if_and_8_cse = PECoreRun_wen & and_626_cse;
  assign rva_in_reg_rw_and_12_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & while_stage_0_9;
  assign input_mem_banks_read_read_data_and_27_cse = PECoreRun_wen & and_dcpl_344
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5) & input_read_req_valid_lpi_1_dfm_1_7;
  assign input_mem_banks_read_read_data_and_69_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_70_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_71_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_72_enex5 = input_mem_banks_read_read_data_and_27_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse = PECoreRun_wen & and_dcpl_348
      & and_dcpl_343 & and_dcpl_347;
  assign and_352_cse = PECore_UpdateFSM_switch_lp_equal_tmp_3_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign input_read_req_valid_and_3_cse = PECoreRun_wen & and_dcpl_344;
  assign PECore_DecodeAxiRead_switch_lp_and_15_cse = PECoreRun_wen & (~(rva_in_reg_rw_sva_7
      | rva_in_reg_rw_sva_st_1_7)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & and_dcpl_347;
  assign rva_out_reg_data_and_243_enex5 = rva_out_reg_data_and_89_ssc & reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_244_enex5 = rva_out_reg_data_and_89_ssc & reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  assign weight_port_read_out_data_and_168_cse = PECoreRun_wen & and_dcpl_343 & while_stage_0_9
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  assign weight_port_read_out_data_and_206_enex5 = weight_port_read_out_data_and_168_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_2_enexo;
  assign weight_port_read_out_data_and_207_enex5 = weight_port_read_out_data_and_168_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  assign rva_out_reg_data_and_245_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_246_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_247_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_62_48_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_248_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_255_240_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_249_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_239_224_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_250_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_223_208_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_251_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_207_192_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_252_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_191_176_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_253_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_175_160_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_254_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_159_144_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_255_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_143_128_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_256_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_127_112_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_257_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_111_96_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_258_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_95_80_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_259_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_79_64_sva_dfm_4_2_enexo;
  assign rva_in_reg_rw_and_15_cse = PECoreRun_wen & and_dcpl_367;
  assign input_mem_banks_read_read_data_and_36_cse = PECoreRun_wen & and_dcpl_372
      & input_read_req_valid_lpi_1_dfm_1_6 & while_stage_0_8;
  assign input_mem_banks_read_read_data_and_73_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_74_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_75_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_76_enex5 = input_mem_banks_read_read_data_and_36_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse = PECoreRun_wen & and_dcpl_371
      & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 | rva_in_reg_rw_sva_6))
      & (~ input_read_req_valid_lpi_1_dfm_1_6) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5
      & while_stage_0_8;
  assign input_read_req_valid_and_4_cse = PECoreRun_wen & and_dcpl_371 & while_stage_0_8;
  assign PECore_DecodeAxiRead_switch_lp_and_19_cse = PECoreRun_wen & and_dcpl_372
      & and_dcpl_380 & while_stage_0_8;
  assign rva_out_reg_data_and_108_ssc = PECoreRun_wen & and_dcpl_372 & and_dcpl_380
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_6) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5
      & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6)
      & (~ rva_in_reg_rw_sva_st_6) & while_stage_0_8;
  assign rva_out_reg_data_and_260_enex5 = rva_out_reg_data_and_108_ssc & reg_rva_out_reg_data_30_25_sva_dfm_4_enexo;
  assign rva_out_reg_data_and_261_enex5 = rva_out_reg_data_and_108_ssc & reg_rva_out_reg_data_23_17_sva_dfm_4_enexo;
  assign rva_out_reg_data_and_262_enex5 = rva_out_reg_data_and_108_ssc & reg_rva_out_reg_data_15_9_sva_dfm_6_enexo;
  assign weight_port_read_out_data_and_170_cse = PECoreRun_wen & and_dcpl_371 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4
      & while_stage_0_8;
  assign weight_port_read_out_data_and_208_enex5 = weight_port_read_out_data_and_170_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_263_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_264_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_265_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_62_48_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_266_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_255_240_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_267_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_239_224_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_268_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_223_208_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_269_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_207_192_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_270_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_191_176_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_271_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_175_160_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_272_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_159_144_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_273_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_143_128_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_274_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_127_112_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_275_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_111_96_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_276_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_95_80_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_277_enex5 = input_read_req_valid_and_4_cse & reg_rva_out_reg_data_79_64_sva_dfm_4_1_enexo;
  assign input_mem_banks_read_read_data_and_45_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1
      & and_dcpl_395;
  assign input_mem_banks_read_read_data_and_77_enex5 = input_mem_banks_read_read_data_and_45_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  assign input_mem_banks_read_read_data_and_78_enex5 = input_mem_banks_read_read_data_and_45_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1;
  assign input_mem_banks_read_read_data_and_79_enex5 = input_mem_banks_read_read_data_and_45_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2;
  assign input_mem_banks_read_read_data_and_80_enex5 = input_mem_banks_read_read_data_and_45_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse = PECoreRun_wen & while_and_21_cse
      & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4
      & while_stage_0_7 & (~ rva_in_reg_rw_sva_st_1_5);
  assign input_read_req_valid_and_5_cse = PECoreRun_wen & and_dcpl_195 & (~ rva_in_reg_rw_sva_st_1_5);
  assign PECore_DecodeAxiRead_switch_lp_and_23_cse = PECoreRun_wen & and_dcpl_408
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1) & while_stage_0_7
      & (~ rva_in_reg_rw_sva_st_1_5);
  assign rva_out_reg_data_and_128_cse = PECoreRun_wen & and_dcpl_408 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_5)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5
      | rva_in_reg_rw_sva_st_5)) & and_dcpl_395;
  assign rva_out_reg_data_and_278_enex5 = rva_out_reg_data_and_128_cse & reg_rva_out_reg_data_23_17_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_279_enex5 = rva_out_reg_data_and_128_cse & reg_rva_out_reg_data_15_9_sva_dfm_5_enexo;
  assign and_1344_cse = (~(((~((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      | rva_in_reg_rw_sva_6 | (~ while_stage_0_8) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)) | rva_in_reg_rw_sva_st_1_5)
      & rva_in_reg_rw_sva_5)) & weight_mem_run_3_for_aelse_and_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign mux_55_nl = MUX_s_1_2_2(and_dcpl_284, or_tmp, rva_in_reg_rw_sva_st_1_5);
  assign rva_out_reg_data_and_134_cse = PECoreRun_wen & (~ mux_55_nl) & while_stage_0_7;
  assign or_666_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      | rva_in_reg_rw_sva_5;
  assign or_671_nl = while_stage_0_6 | mux_402_cse;
  assign mux_59_nl = MUX_s_1_2_2(mux_402_cse, rva_in_reg_rw_sva_4, while_stage_0_6);
  assign mux_60_nl = MUX_s_1_2_2(or_671_nl, mux_59_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_61_nl = MUX_s_1_2_2(mux_60_nl, or_666_cse, while_stage_0_7);
  assign rva_out_reg_data_and_146_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & mux_61_nl;
  assign nand_83_cse = ~(rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse);
  assign or_1369_nl = rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | nand_83_cse;
  assign or_1368_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign mux_400_nl = MUX_s_1_2_2(or_1369_nl, or_1368_nl, while_stage_0_3);
  assign or_1367_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | reg_rva_in_reg_rw_sva_2_cse;
  assign mux_401_nl = MUX_s_1_2_2(mux_400_nl, or_1367_nl, while_stage_0_4);
  assign or_1366_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | rva_in_reg_rw_sva_3;
  assign mux_402_cse = MUX_s_1_2_2(mux_401_nl, or_1366_nl, while_stage_0_5);
  assign or_1365_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | rva_in_reg_rw_sva_4;
  assign mux_403_cse = MUX_s_1_2_2(mux_402_cse, or_1365_nl, while_stage_0_6);
  assign mux_404_nl = MUX_s_1_2_2(mux_403_cse, or_666_cse, while_stage_0_7);
  assign and_1357_cse = mux_404_nl & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & (~ rva_in_reg_rw_sva_6) & while_stage_0_8 & weight_mem_read_arbxbar_arbiters_next_and_cse;
  assign rva_out_reg_data_and_150_cse = PECoreRun_wen & not_tmp_139 & and_dcpl_423;
  assign rva_out_reg_data_and_280_enex5 = rva_out_reg_data_and_150_cse & reg_rva_out_reg_data_46_40_sva_dfm_1_4_enexo;
  assign rva_out_reg_data_and_281_enex5 = rva_out_reg_data_and_150_cse & reg_rva_out_reg_data_39_36_sva_dfm_1_4_enexo;
  assign and_1372_cse = mux_403_cse & and_dcpl_808 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & PECoreRun_wen & (~ rva_in_reg_rw_sva_5);
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_24_cse = PECoreRun_wen & (~(rva_in_reg_rw_sva_st_1_4
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1)) & (~ rva_in_reg_rw_sva_4)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 & and_dcpl_423;
  assign mux_62_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_6_lpi_1_dfm_1, (~ or_tmp_35),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign PECore_DecodeAxiRead_switch_lp_and_27_cse = PECoreRun_wen & mux_62_nl &
      while_stage_0_6;
  assign rva_out_reg_data_and_166_cse = PECoreRun_wen & not_tmp_139 & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_4)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4)
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 | rva_in_reg_rw_sva_st_4
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)) & and_dcpl_56;
  assign rva_out_reg_data_and_282_enex5 = rva_out_reg_data_and_166_cse & reg_rva_out_reg_data_23_17_sva_dfm_2_enexo;
  assign rva_out_reg_data_and_283_enex5 = rva_out_reg_data_and_166_cse & reg_rva_out_reg_data_15_9_sva_dfm_4_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_28_cse = PECoreRun_wen & and_dcpl_444
      & (~(rva_in_reg_rw_sva_3 | input_read_req_valid_lpi_1_dfm_1_3)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_762_nl = (Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp) & PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign or_674_nl = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp;
  assign mux_63_nl = MUX_s_1_2_2(and_762_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      or_674_nl);
  assign mux_64_nl = MUX_s_1_2_2(mux_63_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1_1);
  assign mux_65_nl = MUX_s_1_2_2(mux_64_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp);
  assign mux_66_nl = MUX_s_1_2_2(mux_65_nl, (~ or_tmp_68), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_29_cse = PECoreRun_wen & mux_66_nl
      & while_stage_0_5;
  assign input_mem_banks_read_read_data_and_55_enex5 = PECoreRun_wen & and_dcpl_444
      & input_read_req_valid_lpi_1_dfm_1_3 & and_dcpl_76 & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo;
  assign mux_67_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, (~ or_tmp_68),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign PECore_DecodeAxiRead_switch_lp_and_31_cse = PECoreRun_wen & mux_67_nl &
      while_stage_0_5;
  assign rva_out_reg_data_and_169_cse = PECoreRun_wen & and_dcpl_457 & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_3
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3))
      & (~(input_read_req_valid_lpi_1_dfm_1_3 | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1))
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 & and_dcpl_76;
  assign rva_out_reg_data_and_284_enex5 = rva_out_reg_data_and_169_cse & reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_285_enex5 = rva_out_reg_data_and_169_cse & reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_172_cse = PECoreRun_wen & and_dcpl_457 & (~ input_read_req_valid_lpi_1_dfm_1_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign rva_out_reg_data_and_286_enex5 = rva_out_reg_data_and_172_cse & reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_287_enex5 = rva_out_reg_data_and_172_cse & reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_288_enex5 = rva_out_reg_data_and_172_cse & reg_rva_out_reg_data_62_48_sva_dfm_1_3_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_33_cse = PECoreRun_wen & and_dcpl_468
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 & and_dcpl_133;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse = PECoreRun_wen & and_dcpl_468
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign input_mem_banks_read_read_data_and_56_enex5 = PECoreRun_wen & or_dcpl_606
      & (~ reg_rva_in_reg_rw_sva_2_cse) & input_read_req_valid_lpi_1_dfm_1_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1;
  assign rva_out_reg_data_and_175_cse = PECoreRun_wen & (~(input_read_req_valid_lpi_1_dfm_1_2
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_2)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2))
      & and_dcpl_133 & (~ reg_rva_in_reg_rw_sva_2_cse);
  assign rva_out_reg_data_and_289_enex5 = rva_out_reg_data_and_175_cse & reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  assign rva_out_reg_data_and_290_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_291_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_292_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_293_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse
      & reg_rva_out_reg_data_62_48_sva_dfm_1_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse = PECoreRun_wen & mux_tmp_69
      & and_dcpl_489;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse = PECoreRun_wen & and_dcpl_489;
  assign rva_out_reg_data_and_182_enex5 = PECoreRun_wen & (~(input_read_req_valid_lpi_1_dfm_1_1
      | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[0])))
      & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[3:1]==3'b010)
      & and_dcpl_495 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_294_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_295_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_296_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_297_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse
      & reg_pe_manager_base_input_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse = PECoreRun_wen & mux_tmp_69
      & and_dcpl_488 & (~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1) &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_46_cse = PECoreRun_wen & and_dcpl_187
      & and_dcpl_189 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_48_cse = PECoreRun_wen & and_dcpl_282
      & (~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])))
      & nand_35_cse;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_52_cse = PECoreRun_wen & (or_dcpl_121
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]!=2'b10)) & and_dcpl_226;
  assign PECore_DecodeAxiRead_switch_lp_mux_21_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[0]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_11,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl
      = PECore_DecodeAxiRead_switch_lp_mux_21_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_34_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_19_nl,
      rva_out_reg_data_0_sva_dfm_6, rva_in_reg_rw_sva_11);
  assign PECore_PushAxiRsp_if_else_mux_27_nl = MUX_s_1_2_2(rva_out_reg_data_mux_34_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_6,
      input_read_req_valid_lpi_1_dfm_1_11);
  assign rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_0_mx0 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_27_nl,
      (weight_port_read_out_data_0_0_sva_dfm_6[0]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl
      = (SC_SRAM_CONFIG[7:1]) & (signext_7_1(~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10))
      & ({{6{PECore_DecodeAxiRead_switch_lp_nor_9_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1});
  assign rva_out_reg_data_7_1_sva_dfm_7 = MUX1HOT_v_7_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl,
      rva_out_reg_data_7_1_sva_dfm_6, input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_6,
      (weight_port_read_out_data_0_0_sva_dfm_6[7:1]), {PECore_PushAxiRsp_if_asn_83
      , PECore_PushAxiRsp_if_asn_85 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9});
  assign PECore_DecodeAxiRead_switch_lp_mux_22_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[8]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_11,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl
      = PECore_DecodeAxiRead_switch_lp_mux_22_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_35_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl,
      rva_out_reg_data_8_sva_dfm_6, rva_in_reg_rw_sva_11);
  assign PECore_PushAxiRsp_if_else_mux_28_nl = MUX_s_1_2_2(rva_out_reg_data_mux_35_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_6,
      input_read_req_valid_lpi_1_dfm_1_11);
  assign rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_8_mx0 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_28_nl,
      (weight_port_read_out_data_0_0_sva_dfm_6[8]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9);
  assign PECore_DecodeAxiRead_switch_lp_mux_18_nl = MUX_v_7_2_2((SC_SRAM_CONFIG[15:9]),
      rva_out_reg_data_15_9_sva_dfm_11, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl
      = MUX_v_7_2_2(7'b0000000, PECore_DecodeAxiRead_switch_lp_mux_18_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign rva_out_reg_data_15_9_sva_dfm_7 = MUX1HOT_v_7_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl,
      rva_out_reg_data_15_9_sva_dfm_6, input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_6,
      (weight_port_read_out_data_0_0_sva_dfm_6[15:9]), {PECore_PushAxiRsp_if_asn_83
      , PECore_PushAxiRsp_if_asn_85 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9});
  assign PECore_DecodeAxiRead_switch_lp_mux_23_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[16]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_9,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl
      = PECore_DecodeAxiRead_switch_lp_mux_23_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_36_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl,
      rva_out_reg_data_16_sva_dfm_6, rva_in_reg_rw_sva_11);
  assign PECore_PushAxiRsp_if_else_mux_29_nl = MUX_s_1_2_2(rva_out_reg_data_mux_36_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_6,
      input_read_req_valid_lpi_1_dfm_1_11);
  assign rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_16_mx0 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_29_nl,
      (reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd_1[0]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9);
  assign PECore_DecodeAxiRead_switch_lp_mux_19_nl = MUX_v_7_2_2((SC_SRAM_CONFIG[23:17]),
      rva_out_reg_data_23_17_sva_dfm_9, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl
      = MUX_v_7_2_2(7'b0000000, PECore_DecodeAxiRead_switch_lp_mux_19_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign rva_out_reg_data_23_17_sva_dfm_7 = MUX1HOT_v_7_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl,
      rva_out_reg_data_23_17_sva_dfm_6, input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_6,
      (reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd_1[7:1]), {PECore_PushAxiRsp_if_asn_83
      , PECore_PushAxiRsp_if_asn_85 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9});
  assign PECore_DecodeAxiRead_switch_lp_mux_24_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[24]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_9,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl
      = PECore_DecodeAxiRead_switch_lp_mux_24_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_38_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl,
      rva_out_reg_data_24_sva_dfm_6, rva_in_reg_rw_sva_11);
  assign PECore_PushAxiRsp_if_else_mux_30_nl = MUX_s_1_2_2(rva_out_reg_data_mux_38_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_6,
      input_read_req_valid_lpi_1_dfm_1_11);
  assign rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_24_mx0 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_30_nl,
      (reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd_1[8]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9);
  assign PECore_DecodeAxiRead_switch_lp_mux_20_nl = MUX_v_4_2_2((SC_SRAM_CONFIG[30:27]),
      rva_out_reg_data_30_25_sva_dfm_9_5_2, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl =
      MUX_v_4_2_2(4'b0000, PECore_DecodeAxiRead_switch_lp_mux_20_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign rva_out_reg_data_30_25_sva_dfm_7_5_2 = MUX1HOT_v_4_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl,
      rva_out_reg_data_30_25_sva_dfm_6_5_2_1, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_6[5:2]),
      (reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd_1[14:11]), {PECore_PushAxiRsp_if_asn_83
      , PECore_PushAxiRsp_if_asn_85 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9});
  assign PECore_DecodeAxiRead_switch_lp_mux_25_nl = MUX_v_2_2_2((SC_SRAM_CONFIG[26:25]),
      rva_out_reg_data_30_25_sva_dfm_9_1_0, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl
      = MUX_v_2_2_2(2'b00, PECore_DecodeAxiRead_switch_lp_mux_25_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign rva_out_reg_data_30_25_sva_dfm_7_1_0 = MUX1HOT_v_2_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl,
      rva_out_reg_data_30_25_sva_dfm_6_1_0_1, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_6[1:0]),
      (reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd_1[10:9]), {PECore_PushAxiRsp_if_asn_83
      , PECore_PushAxiRsp_if_asn_85 , PECore_PushAxiRsp_if_asn_87 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl
      = (SC_SRAM_CONFIG[31]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10)
      & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_37_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl,
      rva_out_reg_data_31_sva_dfm_6, rva_in_reg_rw_sva_11);
  assign PECore_PushAxiRsp_if_else_mux_31_nl = MUX_s_1_2_2(rva_out_reg_data_mux_37_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_6,
      input_read_req_valid_lpi_1_dfm_1_11);
  assign rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_31_mx0 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_31_nl,
      reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9);
  assign PECore_RunScale_and_14_nl = (~ PECore_RunScale_if_for_1_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign PECore_RunScale_and_15_nl = PECore_RunScale_if_for_1_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign act_port_reg_data_31_0_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_31_0_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_23 , PECore_RunScale_and_14_nl , PECore_RunScale_and_15_nl});
  assign PECore_RunScale_and_12_nl = (~ PECore_RunScale_if_for_2_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign PECore_RunScale_and_13_nl = PECore_RunScale_if_for_2_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign act_port_reg_data_63_32_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_63_32_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_23 , PECore_RunScale_and_12_nl , PECore_RunScale_and_13_nl});
  assign PECore_RunScale_and_10_nl = (~ PECore_RunScale_if_for_3_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign PECore_RunScale_and_11_nl = PECore_RunScale_if_for_3_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign act_port_reg_data_95_64_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_95_64_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_23 , PECore_RunScale_and_10_nl , PECore_RunScale_and_11_nl});
  assign PECore_RunScale_and_8_nl = (~ PECore_RunScale_if_for_4_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign PECore_RunScale_and_9_nl = PECore_RunScale_if_for_4_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign act_port_reg_data_127_96_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_127_96_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_23 , PECore_RunScale_and_8_nl , PECore_RunScale_and_9_nl});
  assign PECore_RunScale_and_6_nl = (~ PECore_RunScale_if_for_5_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign PECore_RunScale_and_7_nl = PECore_RunScale_if_for_5_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign act_port_reg_data_159_128_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_159_128_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_23 , PECore_RunScale_and_6_nl , PECore_RunScale_and_7_nl});
  assign PECore_RunScale_and_4_nl = (~ PECore_RunScale_if_for_6_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign PECore_RunScale_and_5_nl = PECore_RunScale_if_for_6_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign act_port_reg_data_191_160_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_191_160_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_23 , PECore_RunScale_and_4_nl , PECore_RunScale_and_5_nl});
  assign PECore_RunScale_and_2_nl = (~ PECore_RunScale_if_for_7_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign PECore_RunScale_and_3_nl = PECore_RunScale_if_for_7_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_11 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_11);
  assign act_port_reg_data_223_192_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_223_192_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_asn_23 , PECore_RunScale_and_2_nl , PECore_RunScale_and_3_nl});
  assign and_537_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_5 & while_stage_0_7;
  assign and_542_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9)
      & while_stage_0_11;
  assign and_572_cse = while_stage_0_13 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11
      & (~ rva_in_reg_rw_sva_st_1_11);
  assign and_576_cse = while_stage_0_13 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11)
      & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_11;
  assign PECore_RunMac_or_nl = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_10)
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_10;
  assign PECore_RunScale_and_nl = (~ PECore_RunScale_if_for_8_operator_32_true_slc_32_1_svs_1)
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_10);
  assign PECore_RunScale_and_1_nl = PECore_RunScale_if_for_8_operator_32_true_slc_32_1_svs_1
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_10 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_10);
  assign act_port_reg_data_255_224_sva_dfm_3 = MUX1HOT_v_32_3_2(act_port_reg_data_255_224_sva,
      (PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_z[42:11]), 32'b10000000000000000000000000000001,
      {PECore_RunMac_or_nl , PECore_RunScale_and_nl , PECore_RunScale_and_1_nl});
  assign weight_port_read_out_data_0_0_sva_dfm_1_mx0w0 = MUX1HOT_v_16_9_2(weight_port_read_out_data_0_0_sva_dfm_2,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , and_1441_cse , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , reg_weight_mem_run_3_for_5_and_148_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_151_itm_2 , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign and_1038_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_3_cse & (~
      or_dcpl_720);
  assign and_1039_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      & (~ or_dcpl_720);
  assign and_1040_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1
      & (~ or_dcpl_720);
  assign and_1041_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_231_itm_1
      & (~ or_dcpl_720);
  assign and_1042_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1
      & (~ or_dcpl_720);
  assign nor_473_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl_720);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 & (~ or_dcpl_720);
  assign mux1h_nl = MUX1HOT_v_16_7_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1,
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1,
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[15:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[15:0]),
      weight_port_read_out_data_0_0_sva_dfm_2, {crossbar_spec_PE_Weight_WordType_8U_8U_for_and_nl
      , and_1038_cse , and_1039_cse , and_1040_cse , and_1041_cse , and_1042_cse
      , nor_473_cse});
  assign not_2443_nl = ~ or_dcpl_720;
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w1 = MUX_v_16_2_2(16'b0000000000000000,
      mux1h_nl, not_2443_nl);
  assign PECore_PushAxiRsp_if_else_mux_26_mx0w2 = MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_278_itm_1 = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign Arbiter_8U_Roundrobin_pick_nand_36_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1)
      & and_dcpl_85)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_26_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1
      & and_dcpl_85;
  assign weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_36_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_36_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_36_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_36_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_36_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_36_cse , Arbiter_8U_Roundrobin_pick_and_26_cse});
  assign weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_85);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign Arbiter_8U_Roundrobin_pick_nand_24_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)
      & and_dcpl_85)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_20_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1
      & and_dcpl_85;
  assign weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_24_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_24_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_24_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_24_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_24_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_24_cse , Arbiter_8U_Roundrobin_pick_and_20_cse});
  assign weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_85);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign Arbiter_8U_Roundrobin_pick_nand_12_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1)
      & and_dcpl_85)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_14_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1
      & and_dcpl_85;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_69_nl = weight_mem_read_arbxbar_arbiters_next_5_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_69_nl,
      weight_mem_read_arbxbar_arbiters_next_5_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_12_cse , Arbiter_8U_Roundrobin_pick_and_14_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl = weight_mem_read_arbxbar_arbiters_next_5_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl,
      weight_mem_read_arbxbar_arbiters_next_5_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_12_cse , Arbiter_8U_Roundrobin_pick_and_14_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl = weight_mem_read_arbxbar_arbiters_next_5_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl,
      weight_mem_read_arbxbar_arbiters_next_5_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_12_cse , Arbiter_8U_Roundrobin_pick_and_14_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_nl = weight_mem_read_arbxbar_arbiters_next_5_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_nl,
      weight_mem_read_arbxbar_arbiters_next_5_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_12_cse , Arbiter_8U_Roundrobin_pick_and_14_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_73_nl = weight_mem_read_arbxbar_arbiters_next_5_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_73_nl,
      weight_mem_read_arbxbar_arbiters_next_5_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_12_cse , Arbiter_8U_Roundrobin_pick_and_14_cse});
  assign weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_85);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign Arbiter_8U_Roundrobin_pick_nand_10_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1)
      & and_dcpl_85)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_13_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1
      & and_dcpl_85;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_nl = weight_mem_read_arbxbar_arbiters_next_4_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_nl,
      weight_mem_read_arbxbar_arbiters_next_4_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_77_nl = weight_mem_read_arbxbar_arbiters_next_4_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_77_nl,
      weight_mem_read_arbxbar_arbiters_next_4_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_nl = weight_mem_read_arbxbar_arbiters_next_4_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_nl,
      weight_mem_read_arbxbar_arbiters_next_4_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_10_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_85);
  assign Arbiter_8U_Roundrobin_pick_nand_55_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1)
      & and_dcpl_85)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_44_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1
      & and_dcpl_85;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_81_nl = weight_mem_read_arbxbar_arbiters_next_3_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_81_nl,
      weight_mem_read_arbxbar_arbiters_next_3_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_55_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_82_cse = weight_mem_read_arbxbar_arbiters_next_3_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_82_cse,
      weight_mem_read_arbxbar_arbiters_next_3_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_55_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_55_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_55_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_85_nl = weight_mem_read_arbxbar_arbiters_next_3_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_85_nl,
      weight_mem_read_arbxbar_arbiters_next_3_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_55_cse , Arbiter_8U_Roundrobin_pick_and_44_cse});
  assign weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_85);
  assign Arbiter_8U_Roundrobin_pick_nand_63_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1)
      & and_dcpl_85)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_52_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1
      & and_dcpl_85;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl = weight_mem_read_arbxbar_arbiters_next_2_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl,
      weight_mem_read_arbxbar_arbiters_next_2_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_63_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl = weight_mem_read_arbxbar_arbiters_next_2_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl,
      weight_mem_read_arbxbar_arbiters_next_2_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_63_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl = weight_mem_read_arbxbar_arbiters_next_2_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl,
      weight_mem_read_arbxbar_arbiters_next_2_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_63_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl = weight_mem_read_arbxbar_arbiters_next_2_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl,
      weight_mem_read_arbxbar_arbiters_next_2_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_63_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl,
      weight_mem_read_arbxbar_arbiters_next_2_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_63_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl = weight_mem_read_arbxbar_arbiters_next_2_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl,
      weight_mem_read_arbxbar_arbiters_next_2_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_63_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_85);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign Arbiter_8U_Roundrobin_pick_nand_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1)
      & and_dcpl_85)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_8_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1
      & and_dcpl_85;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl = weight_mem_read_arbxbar_arbiters_next_1_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl,
      weight_mem_read_arbxbar_arbiters_next_1_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_8_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl = weight_mem_read_arbxbar_arbiters_next_1_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl,
      weight_mem_read_arbxbar_arbiters_next_1_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_8_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_95_nl = weight_mem_read_arbxbar_arbiters_next_1_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_95_nl,
      weight_mem_read_arbxbar_arbiters_next_1_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_8_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl,
      weight_mem_read_arbxbar_arbiters_next_1_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_8_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_nl,
      weight_mem_read_arbxbar_arbiters_next_1_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_8_cse});
  assign weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_85);
  assign Arbiter_8U_Roundrobin_pick_nand_85_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1)
      & and_dcpl_85)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_74_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1
      & and_dcpl_85;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_98_nl = weight_mem_read_arbxbar_arbiters_next_0_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_98_nl,
      weight_mem_read_arbxbar_arbiters_next_0_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_85_cse , Arbiter_8U_Roundrobin_pick_and_74_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_99_nl = weight_mem_read_arbxbar_arbiters_next_0_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_99_nl,
      weight_mem_read_arbxbar_arbiters_next_0_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_85_cse , Arbiter_8U_Roundrobin_pick_and_74_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl = weight_mem_read_arbxbar_arbiters_next_0_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl,
      weight_mem_read_arbxbar_arbiters_next_0_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_85_cse , Arbiter_8U_Roundrobin_pick_and_74_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl = weight_mem_read_arbxbar_arbiters_next_0_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl,
      weight_mem_read_arbxbar_arbiters_next_0_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_85_cse , Arbiter_8U_Roundrobin_pick_and_74_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl = weight_mem_read_arbxbar_arbiters_next_0_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_102_nl,
      weight_mem_read_arbxbar_arbiters_next_0_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_85_cse , Arbiter_8U_Roundrobin_pick_and_74_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_103_nl = weight_mem_read_arbxbar_arbiters_next_0_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_103_nl,
      weight_mem_read_arbxbar_arbiters_next_0_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1,
      {and_dcpl_76 , Arbiter_8U_Roundrobin_pick_nand_85_cse , Arbiter_8U_Roundrobin_pick_and_74_cse});
  assign weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_85);
  assign pe_manager_base_weight_sva_mx1_3_0 = MUX_v_4_2_2((pe_manager_base_weight_sva[3:0]),
      (pe_manager_base_weight_sva_dfm_3_1[3:0]), while_stage_0_5);
  assign pe_manager_base_weight_sva_mx2 = MUX_v_15_2_2(pe_manager_base_weight_sva,
      pe_manager_base_weight_sva_dfm_3_1, while_stage_0_5);
  assign pe_manager_base_weight_sva_mx3_0 = MUX_s_1_2_2((pe_manager_base_weight_sva[0]),
      (pe_manager_base_weight_sva_dfm_3_1[0]), while_stage_0_5);
  assign nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000001;
  assign PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_1_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000001;
  assign operator_15_false_acc_nl = nl_operator_15_false_acc_nl[13:0];
  assign weight_read_addrs_2_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000011;
  assign PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_3_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_1_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:2])}) + 13'b0000000000001;
  assign operator_15_false_acc_1_nl = nl_operator_15_false_acc_1_nl[12:0];
  assign weight_read_addrs_4_14_2_lpi_1_dfm_1_1 = MUX_v_13_2_2(13'b0000000000000,
      operator_15_false_acc_1_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000101;
  assign PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_5_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_2_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000011;
  assign operator_15_false_acc_2_nl = nl_operator_15_false_acc_2_nl[13:0];
  assign weight_read_addrs_6_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_2_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000111;
  assign PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_7_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112, and_dcpl_588);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97, and_115_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign and_665_nl = (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5])));
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82, and_665_nl);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl
      & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_5_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_5_tmp = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67, and_122_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign and_658_nl = (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])));
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52, and_658_nl);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl
      & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign and_651_nl = (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])))
      & and_dcpl_635;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37, and_651_nl);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl
      & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign and_644_nl = (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])));
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22, and_644_nl);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl
      & or_185_cse;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_30_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign and_637_nl = (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])))
      & and_dcpl_621;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7, and_637_nl);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl
      & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1 = (state_2_1_sva[0]) & (~((state_2_1_sva[1])
      | state_0_sva));
  assign state_mux_1_cse = MUX_v_2_2_2(state_2_1_sva, state_2_1_sva_dfm_1, while_stage_0_3);
  assign state_0_sva_mx1 = MUX_s_1_2_2(PECore_UpdateFSM_next_state_0_lpi_1_dfm_4,
      state_0_sva, or_dcpl_637);
  assign pe_config_manager_counter_sva_mx1 = MUX_v_4_2_2(pe_config_manager_counter_sva,
      pe_config_manager_counter_sva_dfm_3_1, and_1227_cse);
  assign PECore_PushOutput_PECore_PushOutput_if_and_svs_1 = (state_mux_1_cse[1])
      & (~((state_mux_1_cse[0]) | state_0_sva_mx1));
  assign PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1 = ~(PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_142_cse);
  assign pe_config_input_counter_and_cse = while_if_and_tmp_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign nl_operator_8_false_acc_nl = pe_config_input_counter_sva + 8'b00000001;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[7:0];
  assign pe_config_UpdateInputCounter_not_nl = ~ pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl = MUX_v_8_2_2(8'b00000000,
      operator_8_false_acc_nl, pe_config_UpdateInputCounter_not_nl);
  assign pe_config_input_counter_nand_nl = ~(while_stage_0_3 & (~((~(PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1285_cse_1)));
  assign pe_config_input_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_input_counter_sva,
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl, pe_config_input_counter_sva_dfm_1,
      {pe_config_input_counter_nand_nl , and_352_cse , pe_config_input_counter_and_cse});
  assign nl_operator_8_false_1_acc_nl = pe_config_output_counter_sva + 8'b00000001;
  assign operator_8_false_1_acc_nl = nl_operator_8_false_1_acc_nl[7:0];
  assign pe_config_UpdateManagerCounter_if_not_9_nl = ~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl
      = MUX_v_8_2_2(8'b00000000, operator_8_false_1_acc_nl, pe_config_UpdateManagerCounter_if_not_9_nl);
  assign pe_config_output_counter_nand_nl = ~(while_stage_0_3 & (~((~(and_1437_cse
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1285_cse_1)));
  assign while_and_164_nl = and_1437_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign pe_config_output_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_output_counter_sva,
      pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl,
      pe_config_output_counter_sva_dfm_1, {pe_config_output_counter_nand_nl , while_and_164_nl
      , pe_config_input_counter_and_cse});
  assign and_626_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_if_and_2_m1c = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & and_626_cse;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl
      = pe_config_is_zero_first_sva & (~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1);
  assign while_if_or_nl = (~((~((~ PECore_UpdateFSM_switch_lp_equal_tmp_5_1) & and_626_cse))
      & while_stage_0_3)) | ((~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1)
      & while_if_and_2_m1c);
  assign while_if_and_4_nl = pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
      & while_if_and_2_m1c;
  assign pe_config_is_zero_first_sva_mx1 = MUX1HOT_s_1_3_2(while_if_mux_27_itm_1,
      pe_config_is_zero_first_sva, pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl,
      {and_dcpl_172 , while_if_or_nl , while_if_and_4_nl});
  assign PECore_UpdateFSM_switch_lp_equal_tmp_6 = state_0_sva_mx1 & (state_mux_1_cse==2'b00);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1 = (state_mux_1_cse[0])
      & (~((state_mux_1_cse[1]) | state_0_sva_mx1));
  assign pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1
      = ~((pe_config_manager_counter_sva_mx1 != (operator_4_false_acc_sdt_sva_1[3:0]))
      | (operator_4_false_acc_sdt_sva_1[4]));
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0110);
  assign weight_port_read_out_data_0_3_sva_mx0 = MUX1HOT_v_16_3_2(weight_port_read_out_data_0_3_sva_dfm_1,
      weight_port_read_out_data_0_3_sva_dfm_1_1, weight_port_read_out_data_0_3_sva,
      {and_dcpl_367 , and_dcpl_320 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_2_sva_mx0 = MUX1HOT_v_16_3_2(weight_port_read_out_data_0_2_sva_dfm_1,
      weight_port_read_out_data_0_2_sva_dfm_1_1, weight_port_read_out_data_0_2_sva,
      {and_dcpl_367 , and_dcpl_320 , (~ while_stage_0_8)});
  assign mux1h_5_nl = MUX1HOT_v_16_7_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[63:48]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63:48]),
      weight_port_read_out_data_0_3_sva_mx0, {and_1017_cse , and_1018_cse , and_1019_cse
      , and_1020_cse , and_1021_cse , and_1022_cse , nor_472_cse});
  assign not_2445_nl = ~ or_dcpl;
  assign weight_port_read_out_data_0_3_sva_dfm_2 = MUX_v_16_2_2(16'b0000000000000000,
      mux1h_5_nl, not_2445_nl);
  assign and_1053_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_28 & (~ or_dcpl_720);
  assign mux1h_6_nl = MUX1HOT_v_16_7_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[47:32]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[47:32]),
      weight_port_read_out_data_0_2_sva_mx0, {and_1053_nl , and_1038_cse , and_1039_cse
      , and_1040_cse , and_1041_cse , and_1042_cse , nor_473_cse});
  assign not_2447_nl = ~ or_dcpl_720;
  assign weight_port_read_out_data_0_2_sva_dfm_2 = MUX_v_16_2_2(16'b0000000000000000,
      mux1h_6_nl, not_2447_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2!=3'b000));
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  assign weight_mem_run_3_for_land_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1);
  assign weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6,
      or_dcpl_636);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0,
      or_dcpl_636);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5,
      or_dcpl_636);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1,
      or_dcpl_636);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4,
      or_dcpl_636);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2,
      or_dcpl_636);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3,
      or_dcpl_636);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_1_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0101);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1 = (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp;
  assign weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & weight_mem_read_arbxbar_xbar_1_for_3_8_for_4_or_cse;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  assign weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b111)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b100)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_40_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b011)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b010)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b001)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_mx0w0 = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_359_itm_1
      & (pe_manager_base_weight_sva[1:0]==2'b10) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign weight_mem_run_3_for_land_1_lpi_1_dfm_1_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1 = MUX_v_3_2_2(3'b000,
      (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0]), weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp = MUX_s_1_8_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp
      | (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp));
  assign while_and_234_rgt = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_238_rgt = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_242_rgt = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_246_rgt = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_250_rgt = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_254_rgt = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_258_rgt = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_262_rgt = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_266_rgt = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_270_rgt = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_274_rgt = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_278_rgt = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_282_rgt = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_286_rgt = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_290_rgt = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_294_rgt = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_298_rgt = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_302_rgt = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_306_rgt = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_310_rgt = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_314_rgt = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_318_rgt = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_322_rgt = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_326_rgt = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_330_rgt = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_334_rgt = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_338_rgt = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_342_rgt = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_346_rgt = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_350_rgt = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_354_rgt = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_358_rgt = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_362_rgt = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_366_rgt = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_370_rgt = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_374_rgt = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_378_rgt = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_382_rgt = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_386_rgt = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_390_rgt = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_394_rgt = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_398_rgt = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_402_rgt = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_406_rgt = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_410_rgt = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_414_rgt = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_418_rgt = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_422_rgt = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_426_rgt = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_430_rgt = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_434_rgt = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_438_rgt = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_442_rgt = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_446_rgt = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_450_rgt = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_454_rgt = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_458_rgt = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_462_rgt = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_466_rgt = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_470_rgt = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_474_rgt = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_478_rgt = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_482_rgt = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_486_rgt = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_490_rgt = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_494_rgt = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_498_rgt = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_502_rgt = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_506_rgt = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_510_rgt = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_514_rgt = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_518_rgt = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_522_rgt = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_526_rgt = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_530_rgt = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_534_rgt = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_538_rgt = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_542_rgt = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_546_rgt = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_550_rgt = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_554_rgt = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_558_rgt = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_562_rgt = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_566_rgt = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_570_rgt = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_574_rgt = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_578_rgt = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_582_rgt = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_586_rgt = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_590_rgt = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_594_rgt = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_598_rgt = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_602_rgt = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_606_rgt = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_610_rgt = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_614_rgt = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_618_rgt = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_622_rgt = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_626_rgt = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_630_rgt = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 &
      (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_634_rgt = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_638_rgt = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_642_rgt = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_646_rgt = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_650_rgt = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_654_rgt = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_658_rgt = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_662_rgt = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_666_rgt = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_670_rgt = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_674_rgt = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_678_rgt = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_682_rgt = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_686_rgt = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_690_rgt = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_694_rgt = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_698_rgt = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_702_rgt = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_706_rgt = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_710_rgt = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_714_rgt = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_718_rgt = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_722_rgt = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_726_rgt = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_730_rgt = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_734_rgt = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_738_rgt = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_742_rgt = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_746_rgt = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_750_rgt = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_754_rgt = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_758_rgt = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_762_rgt = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_766_rgt = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_770_rgt = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_774_rgt = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_778_rgt = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_782_rgt = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_786_rgt = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_790_rgt = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_794_rgt = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_798_rgt = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_802_rgt = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_806_rgt = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_810_rgt = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_814_rgt = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_818_rgt = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_822_rgt = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_826_rgt = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_830_rgt = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_834_rgt = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_838_rgt = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_842_rgt = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_846_rgt = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_850_rgt = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_854_rgt = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_858_rgt = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_862_rgt = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_866_rgt = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_870_rgt = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_874_rgt = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_878_rgt = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_882_rgt = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_886_rgt = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_890_rgt = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_894_rgt = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_898_rgt = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_902_rgt = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_906_rgt = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_910_rgt = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_914_rgt = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_918_rgt = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_922_rgt = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_926_rgt = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_930_rgt = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_934_rgt = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_938_rgt = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_942_rgt = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_946_rgt = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_950_rgt = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_954_rgt = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_958_rgt = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_962_rgt = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_966_rgt = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_970_rgt = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_974_rgt = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_978_rgt = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_982_rgt = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_986_rgt = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_990_rgt = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_994_rgt = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_998_rgt = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1002_rgt = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1006_rgt = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1010_rgt = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1014_rgt = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1018_rgt = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1022_rgt = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1026_rgt = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1030_rgt = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1034_rgt = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1038_rgt = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1042_rgt = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1046_rgt = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1050_rgt = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1054_rgt = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1058_rgt = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1062_rgt = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1066_rgt = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1070_rgt = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1074_rgt = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1078_rgt = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1082_rgt = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1086_rgt = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1090_rgt = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1094_rgt = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1098_rgt = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1102_rgt = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1106_rgt = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1110_rgt = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1114_rgt = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1118_rgt = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1122_rgt = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1126_rgt = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1130_rgt = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1134_rgt = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1138_rgt = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1142_rgt = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1146_rgt = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1150_rgt = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1154_rgt = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1158_rgt = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1162_rgt = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1166_rgt = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1170_rgt = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1174_rgt = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1178_rgt = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1182_rgt = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1186_rgt = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1190_rgt = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1194_rgt = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1198_rgt = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1202_rgt = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1206_rgt = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1210_rgt = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1214_rgt = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1218_rgt = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1222_rgt = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1226_rgt = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1230_rgt = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1234_rgt = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1238_rgt = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1242_rgt = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1246_rgt = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1250_rgt = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_and_1254_rgt = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign pe_manager_base_input_sva_mx1 = MUX_v_15_2_2(pe_manager_base_input_sva,
      pe_manager_base_input_sva_dfm_3_1, while_stage_0_3);
  assign PECore_PushAxiRsp_mux_27_nl = MUX_s_1_2_2(pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2,
      PECore_PushAxiRsp_mux_10_itm_1, rva_in_reg_rw_sva_5);
  assign PECore_PushAxiRsp_if_else_mux_10_mx0w2 = MUX_s_1_2_2(PECore_PushAxiRsp_mux_27_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1);
  assign while_if_while_if_and_24_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_255_240_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_255_240_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_24_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[255:240]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_239_2000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_25_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_239_224_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_239_224_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_25_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[239:224]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_223_2000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_26_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_223_208_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_223_208_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_26_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[223:208]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_207_1000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_27_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_207_192_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_207_192_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_27_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[207:192]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_191_1000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_28_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_191_176_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_191_176_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_28_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[191:176]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_175_1000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_29_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_175_160_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_175_160_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_29_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[175:160]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_159_1000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_30_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_159_144_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_159_144_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_30_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[159:144]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_143_1000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_31_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_143_128_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_143_128_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_31_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[143:128]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_127_1000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_32_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_127_112_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_127_112_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_32_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_111_9000000,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_33_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_111_96_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_111_96_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_33_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_95_80_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_34_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_95_80_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_95_80_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_34_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_79_64_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign while_if_while_if_and_35_nl = MUX_v_16_2_2(16'b0000000000000000, rva_out_reg_data_79_64_sva_dfm_6,
      rva_in_reg_rw_sva_5);
  assign rva_out_reg_data_79_64_sva_dfm_4_mx0w0 = MUX1HOT_v_16_3_2(while_if_while_if_and_35_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_63_48_sva_1,
      {PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 , PECore_PushAxiRsp_if_asn_91
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
  assign rva_out_reg_data_62_48_sva_dfm_6_mx1 = MUX_v_15_2_2(rva_out_reg_data_62_48_sva_dfm_4_1,
      rva_out_reg_data_62_48_sva_dfm_6, or_dcpl_706);
  assign rva_out_reg_data_46_40_sva_dfm_6_mx1 = MUX_v_7_2_2(rva_out_reg_data_46_40_sva_dfm_4_1,
      rva_out_reg_data_46_40_sva_dfm_6, or_dcpl_706);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1 = MUX_v_4_2_2(rva_out_reg_data_39_36_sva_dfm_4_1,
      rva_out_reg_data_39_36_sva_dfm_6, or_dcpl_706);
  assign PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
      & PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3
      | and_279_cse);
  assign PECore_DecodeAxiRead_switch_lp_nor_tmp_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_RunScale_PECore_RunScale_if_and_1_svs_1 = (state_mux_1_cse[0]) &
      state_0_sva_mx1 & (~ (state_mux_1_cse[1]));
  assign PECore_DecodeAxiRead_switch_lp_nor_9_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_11
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_11 | PECore_DecodeAxiRead_switch_lp_nor_tmp_11);
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1 = ~(input_read_req_valid_lpi_1_dfm_1_11
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9);
  assign PECore_RunScale_if_for_7_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_2_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_6_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_3_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_5_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_4_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_4_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_5_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_3_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_6_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_2_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_7_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign PECore_RunScale_if_for_1_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0 = MUX_v_256_2_2(weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0 = MUX_v_240_2_2(weight_mem_banks_read_1_read_data_lpi_1_dfm_1_255_16,
      (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[255:16]), weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_load_store_1_for_else_else_and_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_or_nl = (weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1);
  assign weight_mem_banks_load_store_1_for_else_else_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9 = MUX1HOT_v_16_6_2(BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1,
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1,
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[15:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[15:0]),
      {weight_mem_banks_load_store_1_for_else_else_and_nl , weight_mem_banks_load_store_1_for_else_else_or_nl
      , weight_mem_banks_load_store_1_for_else_else_and_4_nl , weight_mem_banks_load_store_1_for_else_else_and_6_nl
      , weight_mem_banks_load_store_1_for_else_else_and_8_nl , weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2});
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1 = (~(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_sva_1 | mux_129_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_sva_1 & (~ mux_129_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_sva_1 | mux_136_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_sva_1 & (~ mux_136_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_sva_1) & and_dcpl_680;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_sva_1 & and_dcpl_680;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]),
      {mux_tmp_126 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_sva_1,
      {mux_tmp_126 , (~ mux_129_itm) , (~ mux_136_itm) , and_dcpl_680});
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  assign mux_145_nl = MUX_s_1_2_2(or_tmp_177, or_tmp_174, while_stage_0_5);
  assign or_887_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva | or_tmp_177;
  assign or_884_nl = while_mux_1472_tmp | or_tmp_174;
  assign mux_144_nl = MUX_s_1_2_2(or_887_nl, or_884_nl, while_stage_0_5);
  assign mux_146_nl = MUX_s_1_2_2(mux_145_nl, mux_144_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl,
      mux_146_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 | mux_158_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 & (~ mux_158_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 | mux_172_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 & (~ mux_172_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1) & and_dcpl_683;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 & and_dcpl_683;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]),
      {mux_tmp_149 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1,
      {mux_tmp_149 , (~ mux_158_itm) , (~ mux_172_itm) , and_dcpl_683});
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  assign mux_181_nl = MUX_s_1_2_2(or_tmp_224, or_tmp_219, while_stage_0_5);
  assign or_934_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | or_tmp_224;
  assign or_929_nl = while_mux_1465_tmp | or_tmp_219;
  assign mux_180_nl = MUX_s_1_2_2(or_934_nl, or_929_nl, while_stage_0_5);
  assign mux_182_nl = MUX_s_1_2_2(mux_181_nl, mux_180_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl,
      mux_182_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1) & and_dcpl_686;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 & and_dcpl_686;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1) & and_dcpl_690;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 & and_dcpl_690;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1) & and_dcpl_696;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 & and_dcpl_696;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp,
      weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]),
      {or_dcpl_710 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1,
      {or_dcpl_710 , and_dcpl_686 , and_dcpl_690 , and_dcpl_696});
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign and_707_nl = (~ mux_tmp_189) & and_dcpl_689;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl,
      and_707_nl);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      = weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      = weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      = weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1) & and_dcpl_698;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 & and_dcpl_698;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1) & and_dcpl_701;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 & and_dcpl_701;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1) & and_dcpl_707;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 & and_dcpl_707;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp,
      weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]),
      {or_dcpl_711 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1,
      {or_dcpl_711 , and_dcpl_698 , and_dcpl_701 , and_dcpl_707});
  assign and_997_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  assign and_999_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) & while_mux_1451_tmp;
  assign and_996_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  assign and_998_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]) & while_mux_1454_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign nor_464_nl = ~(and_996_cse | and_997_cse | or_tmp_242);
  assign nor_465_nl = ~(and_998_cse | and_999_cse | or_tmp_238);
  assign mux_206_nl = MUX_s_1_2_2(nor_464_nl, nor_465_nl, while_stage_0_5);
  assign and_718_nl = mux_206_nl & and_dcpl_700;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl,
      and_718_nl);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      = weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      = weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | (weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]));
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_24_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1) & and_dcpl_711;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 & and_dcpl_711;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1) & and_dcpl_714;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 & and_dcpl_714;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1) & and_dcpl_721;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 & and_dcpl_721;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp,
      Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1, (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]), {or_dcpl_713 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_24_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_26_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1,
      operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1, {or_dcpl_713 , and_dcpl_711
      , and_dcpl_714 , and_dcpl_721});
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | (weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign or_1010_nl = weight_mem_read_arbxbar_arbiters_next_3_5_sva | or_tmp_294;
  assign or_1009_nl = while_mux_1445_tmp | mux_tmp_237;
  assign mux_239_nl = MUX_s_1_2_2(or_1010_nl, or_1009_nl, while_stage_0_5);
  assign mux_240_nl = MUX_s_1_2_2(mux_tmp_238, mux_239_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign and_732_nl = (~ mux_240_nl) & and_dcpl_713;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl,
      and_732_nl);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 | mux_257_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 & (~ mux_257_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 | mux_276_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 & (~ mux_276_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1) & and_dcpl_725;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 & and_dcpl_725;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]),
      {mux_tmp_247 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1,
      {mux_tmp_247 , (~ mux_257_itm) , (~ mux_276_itm) , and_dcpl_725});
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1;
  assign mux_286_nl = MUX_s_1_2_2(mux_tmp_266, mux_tmp_264, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_nl,
      mux_286_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1) & and_dcpl_728;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 & and_dcpl_728;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1) & and_dcpl_732;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 & and_dcpl_732;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1) & and_dcpl_738;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 & and_dcpl_738;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp,
      weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]),
      {or_dcpl_715 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1,
      {or_dcpl_715 , and_dcpl_728 , and_dcpl_732 , and_dcpl_738});
  assign and_1000_cse = weight_mem_read_arbxbar_arbiters_next_1_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign and_1001_cse = while_mux_1435_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign nor_466_nl = ~(and_1000_cse | nor_tmp_199);
  assign nor_467_nl = ~(and_1001_cse | nor_tmp_197);
  assign mux_294_nl = MUX_s_1_2_2(nor_466_nl, nor_467_nl, while_stage_0_5);
  assign and_749_nl = mux_294_nl & and_dcpl_731;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl,
      and_749_nl);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      = weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      = weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      = weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 | mux_311_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 & (~ mux_311_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 | mux_324_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 & (~ mux_324_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_46_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1) & and_dcpl_742;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_47_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 & and_dcpl_742;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]),
      {mux_tmp_301 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_46_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_47_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1,
      {mux_tmp_301 , (~ mux_311_itm) , (~ mux_324_itm) , and_dcpl_742});
  assign and_1007_cse = Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign and_1008_cse = Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign and_1009_cse = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign and_1002_cse = Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign and_1004_cse = Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign and_1003_cse = Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]);
  assign and_1006_cse = Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign and_1005_cse = Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign or_1140_cse = and_1003_cse | and_1004_cse | and_1005_cse | and_1006_cse
      | and_1007_cse | and_1008_cse;
  assign mux_335_cse = MUX_s_1_2_2(or_tmp_377, or_1140_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1;
  assign or_1141_nl = and_1002_cse | mux_335_cse;
  assign or_1129_nl = and_1009_cse | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign mux_334_nl = MUX_s_1_2_2(or_tmp_418, or_1129_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign mux_336_nl = MUX_s_1_2_2(or_1141_nl, mux_334_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_337_nl = MUX_s_1_2_2(or_tmp_418, mux_336_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl,
      mux_337_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_125_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = (pe_manager_base_weight_sva_mx2[14:4])
      + PEManager_15U_GetWeightAddr_else_acc_3_1;
  assign PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1[10:0];
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_1_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_1_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_1_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_1_sva_1 | (weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 | (weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 | (weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]));
  assign operator_7_false_1_operator_7_false_1_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 | (weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]));
  assign weight_read_addrs_0_3_0_lpi_1_dfm_4 = MUX_v_4_2_2(4'b0000, pe_manager_base_weight_sva_mx1_3_0,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_4_false_acc_sdt_sva_1 = conv_u2s_4_5(pe_config_num_manager_sva)
      + 5'b11111;
  assign operator_4_false_acc_sdt_sva_1 = nl_operator_4_false_acc_sdt_sva_1[4:0];
  assign while_and_1285_cse_1 = (~ while_if_and_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_if_and_tmp_1 = PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      = ~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl = start_PopNB_mioi_data_rsc_z_mxwt
      & pe_config_is_valid_sva & start_PopNB_mioi_return_rsc_z_mxwt;
  assign PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl = pe_config_is_zero_first_sva
      & pe_manager_zero_active_sva;
  assign PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl = ~(pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign PECore_UpdateFSM_switch_lp_mux1h_15_nl = MUX1HOT_s_1_4_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl,
      PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl, pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1,
      PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl, {PECore_UpdateFSM_switch_lp_and_7_itm_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_2_1 , PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_5_1});
  assign PECore_UpdateFSM_next_state_0_lpi_1_dfm_4 = PECore_UpdateFSM_switch_lp_mux1h_15_nl
      & PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  assign pe_config_UpdateManagerCounter_if_if_unequal_tmp = pe_config_output_counter_sva
      != (operator_8_false_acc_sdt_sva_1[7:0]);
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      = ~(pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]));
  assign input_write_req_valid_lpi_1_dfm_5 = PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      & PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1 = ~(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign PECore_RunScale_if_for_8_operator_32_true_slc_32_1_svs_1 = $signed((PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_1_z[42:11]))
      < $signed(32'b10000000000000000000000000000001);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[255:240]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[255:240]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[239:224]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[255:240]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[255:240]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[239:224]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[255:240]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[255:240]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[239:224]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[239:224]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[239:224]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[223:208]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[223:208]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[223:208]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[207:192]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[207:192]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[207:192]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[191:176]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[191:176]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[191:176]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[175:160]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[175:160]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[175:160]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[159:144]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[159:144]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[159:144]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[143:128]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[143:128]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[143:128]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[127:112]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[111:96]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[95:80]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[79:64]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[63:48]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[47:32]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[31:16]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[15:0]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000
      = MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[63:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126 , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , reg_weight_mem_run_3_for_5_and_148_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[79:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126 , reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_147_itm_2_cse , reg_weight_mem_run_3_for_5_and_148_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_149_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2 , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[95:80]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_148_itm_2_cse , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_69_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[111:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_69_nl
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_148_itm_2_cse , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[143:128]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[143:128]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[127:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_148_itm_2_cse , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[159:144]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[159:144]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[143:128]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_148_itm_2_cse , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[175:160]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[175:160]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[159:144]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2 , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[191:176]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[191:176]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[175:160]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_148_itm_2_cse , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[207:192]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[207:192]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[191:176]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2 , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[223:208]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[223:208]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[207:192]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2 , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[239:224]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[239:224]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[223:208]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_128
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2
      , reg_weight_mem_run_3_for_5_and_152_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[255:240]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[255:240]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[239:224]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_128
      , reg_weight_mem_run_3_for_5_and_146_itm_2_cse , reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_2 , reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_3 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_3
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_3});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[15:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[31:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[47:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[63:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[79:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[95:80]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[111:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_nl , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[143:128]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[143:128]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[127:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[159:144]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[159:144]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[143:128]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[175:160]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[175:160]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[159:144]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[191:176]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[191:176]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[175:160]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[207:192]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[207:192]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[191:176]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[223:208]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[223:208]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[207:192]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[239:224]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[239:224]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[223:208]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse = reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_453
      , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_1_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[15:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_453
      , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_6_itm_1_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[31:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_453
      , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_15_itm_1_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[47:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_453
      , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , reg_weight_mem_run_3_for_5_and_16_itm_1_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[63:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_453
      , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_336_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[79:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse , weight_mem_run_3_for_5_asn_453
      , weight_mem_run_3_for_5_asn_455 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_328_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[95:80]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse
      , weight_mem_run_3_for_5_asn_453 , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_411});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[111:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse
      , weight_mem_run_3_for_5_asn_453 , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_411});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[143:128]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[143:128]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[127:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse
      , weight_mem_run_3_for_5_asn_453 , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , PECore_DecodeAxiRead_switch_lp_nor_tmp_5});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[159:144]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[159:144]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[143:128]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365
      , weight_mem_run_3_for_5_asn_453 , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_411});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[175:160]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[175:160]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[159:144]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse
      , weight_mem_run_3_for_5_asn_453 , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_411});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[191:176]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[191:176]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[175:160]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365
      , weight_mem_run_3_for_5_asn_453 , weight_mem_run_3_for_5_asn_455 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1
      , weight_mem_run_3_for_5_asn_457 , PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5
      , reg_weight_mem_run_3_for_5_and_7_itm_2_cse , PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[207:192]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[207:192]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[191:176]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365
      , weight_mem_run_3_for_5_asn_453 , weight_mem_run_3_for_5_asn_455 , reg_weight_mem_run_3_for_5_and_12_itm_2_cse
      , weight_mem_run_3_for_5_asn_457 , reg_weight_mem_run_3_for_5_and_14_itm_2_cse
      , PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_411});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[223:208]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[223:208]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[207:192]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_361_cse
      , weight_mem_run_3_for_5_asn_453 , weight_mem_run_3_for_5_asn_455 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1
      , weight_mem_run_3_for_5_asn_457 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[15:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[31:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_419});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[47:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_231_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[63:48]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[79:64]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_231_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[95:80]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[111:96]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[143:128]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[143:128]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[143:128]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[127:112]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[159:144]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[159:144]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[159:144]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[143:128]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[175:160]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[175:160]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[175:160]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[159:144]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[191:176]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[191:176]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[191:176]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[175:160]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[207:192]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[207:192]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[207:192]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[191:176]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[223:208]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[223:208]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[223:208]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[207:192]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_419});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014
      = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[239:224]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[239:224]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[239:224]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[223:208]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_419});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b100)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])
      & nor_526_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      | Arbiter_8U_Roundrobin_pick_1_if_1_and_30_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0,
      or_dcpl_717);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      = MUX_s_1_2_2(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0,
      or_dcpl_717);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      = MUX_s_1_2_2(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0,
      or_dcpl_717);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0
      = MUX_s_1_2_2(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0,
      or_dcpl_717);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0,
      or_dcpl_717);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0,
      or_dcpl_717);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0,
      or_dcpl_717);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1 = and_279_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  assign nl_operator_16_false_acc_sdt_sva_1 = conv_u2s_8_9(pe_manager_num_input_sva)
      + 9'b111111111;
  assign operator_16_false_acc_sdt_sva_1 = nl_operator_16_false_acc_sdt_sva_1[8:0];
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1 = ~((state_mux_1_cse!=2'b00)
      | state_0_sva_mx1);
  assign PECore_UpdateFSM_switch_lp_nor_tmp_1 = ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_6 | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1
      | PECore_RunScale_PECore_RunScale_if_and_1_svs_1 | PECore_PushOutput_PECore_PushOutput_if_and_svs_1);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_144_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_111_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[255:240]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_144_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_159_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_127_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[255:240]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_159_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_239_2000000
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_111_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_127_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_145_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_110_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[239:224]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_145_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_160_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_126_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[239:224]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_160_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_223_2000000
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_110_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_126_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_146_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_109_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[223:208]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_146_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_161_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_125_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[223:208]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_161_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_207_1000000
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_109_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_125_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_147_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_108_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[207:192]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_147_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_162_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_124_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[207:192]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_162_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_191_1000000
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_108_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_124_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_148_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_100_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[79:64]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_148_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_163_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_116_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[79:64]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_163_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_63_48_sva_1
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_36_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_68_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_100_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_116_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_149_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_107_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[191:176]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_149_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_164_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_123_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[191:176]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_164_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_175_1000000
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_107_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_123_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_150_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_101_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[95:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_150_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_165_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_117_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[95:80]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_165_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_79_64_sva_1
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_37_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_69_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_101_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_117_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_151_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_106_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[175:160]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_151_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_166_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_122_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[175:160]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_166_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_159_1000000
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_106_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_122_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_152_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_102_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[111:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_152_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_167_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_118_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[111:96]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_167_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_95_80_sva_1
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_102_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_118_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_153_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_105_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[159:144]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_153_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_168_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_121_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[159:144]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_168_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_143_1000000
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_105_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_121_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_154_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_103_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[127:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_154_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_169_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_119_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[127:112]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_169_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_111_9000000
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_39_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_71_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_103_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_119_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_155_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_104_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[143:128]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_155_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_170_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_120_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[143:128]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_170_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_127_1000000
      = MUX_v_16_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_104_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_120_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign while_and_46_tmp = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp
      = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2) | reg_rva_in_reg_rw_sva_2_cse
      | (~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp!=8'b00000000))) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7])));
  assign PECore_DecodeAxiWrite_switch_lp_or_5_cse_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  assign input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_1_0_sva_1 = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]!=2'b00));
  assign input_mem_banks_write_if_for_if_and_stg_1_1_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b01);
  assign input_mem_banks_write_if_for_if_and_stg_1_2_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b10);
  assign input_mem_banks_write_if_for_if_and_stg_1_3_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b11);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign nl_PEManager_15U_GetInputAddr_acc_nl = input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt
      + (pe_manager_base_input_sva[7:0]);
  assign PEManager_15U_GetInputAddr_acc_nl = nl_PEManager_15U_GetInputAddr_acc_nl[7:0];
  assign input_write_addrs_lpi_1_dfm_2 = PEManager_15U_GetInputAddr_acc_nl & ({{7{PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1}},
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1})
      & ({{7{PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1}}, PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1});
  assign input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1 = ~((input_write_addrs_lpi_1_dfm_2[1:0]!=2'b00));
  assign input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b01);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b10);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b11);
  assign PECore_PushAxiRsp_mux_24_nl = MUX_s_1_2_2(PECore_PushAxiRsp_mux_26_itm_1,
      rva_out_reg_data_63_sva_dfm_6, nand_72_cse);
  assign rva_out_reg_data_63_sva_dfm_7 = PECore_PushAxiRsp_mux_24_nl & rva_in_reg_rw_sva_5;
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2
      | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_4 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0011);
  assign PECore_DecodeAxiRead_switch_lp_nor_13_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_not_185 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 =
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:1]!=15'b000000000000000));
  assign PECore_PushAxiRsp_if_asn_83 = (~ rva_in_reg_rw_sva_11) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_85 = rva_in_reg_rw_sva_11 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_87 = input_read_req_valid_lpi_1_dfm_1_11 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9);
  assign PECore_RunMac_asn_23 = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_11)
      | PECore_RunMac_PECore_RunMac_if_and_svs_11;
  assign weight_mem_run_3_for_5_asn_445 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_447 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_449 = (weight_read_addrs_7_lpi_1_dfm_3_2_0[2])
      & nor_500_cse & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_451 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_453 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_455 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_457 = (weight_read_addrs_5_lpi_1_dfm_3_2_0[2])
      & nor_508_cse & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_411 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_419 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign while_and_45_cse = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign while_while_nor_259_cse = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_3 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign while_and_1256_cse = weight_mem_run_3_for_land_1_lpi_1_dfm_3 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign PECore_PushAxiRsp_if_asn_91 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign PECore_PushAxiRsp_if_asn_93 = (~ rva_in_reg_rw_sva_5) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign PECore_PushAxiRsp_if_asn_95 = rva_in_reg_rw_sva_5 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign while_and_21_cse = (~ rva_in_reg_rw_sva_5) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_363 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_14_itm_1
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_365 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_36_itm_1
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_367 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_153 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_157 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_28 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_128 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_3
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_2
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_2
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign Arbiter_8U_Roundrobin_pick_1_mux_583_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1477_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_583_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_584_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1476_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_584_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_585_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1475_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_585_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_586_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1474_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_586_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_587_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1473_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_587_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_588_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1472_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_588_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1471_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_589_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1470_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_589_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_590_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1469_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_590_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_591_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1468_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_591_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_592_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1467_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_592_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_593_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1466_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_593_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_594_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1465_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_594_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1464_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1457_cse_1 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_601_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1456_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_601_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_603_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1454_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_603_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_606_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1451_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_606_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1450_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_611_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1445_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_611_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_619_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1435_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_619_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1429_cse_1 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_dcpl_6 = while_stage_0_12 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_10;
  assign and_dcpl_7 = and_dcpl_6 & (~ rva_in_reg_rw_sva_st_1_10);
  assign and_dcpl_8 = and_dcpl_7 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8
      | rva_in_reg_rw_sva_10 | input_read_req_valid_lpi_1_dfm_1_10));
  assign and_dcpl_24 = while_stage_0_12 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_10);
  assign and_dcpl_40 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & while_stage_0_9;
  assign or_tmp = (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign and_dcpl_45 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7;
  assign and_dcpl_56 = while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign and_dcpl_57 = while_stage_0_6 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_dcpl_76 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_dcpl_85 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_87 = (((Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1) | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1)
      & and_dcpl_85;
  assign and_dcpl_89 = (((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1) | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1)
      & and_dcpl_85;
  assign and_dcpl_91 = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign or_dcpl_32 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse;
  assign and_dcpl_93 = (((or_dcpl_32 | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1) | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1)
      & and_dcpl_85;
  assign and_dcpl_95 = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_97 = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign or_50_cse = ((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1) | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp;
  assign and_dcpl_99 = or_50_cse & and_dcpl_85;
  assign and_dcpl_101 = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign nor_279_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]));
  assign nor_276_cse = ~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]));
  assign nor_280_cse = ~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]));
  assign and_115_cse = nor_280_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]))) & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])));
  assign or_dcpl_47 = (~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_5_tmp)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4);
  assign nor_284_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]));
  assign and_122_cse = nor_284_cse & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])));
  assign or_dcpl_48 = and_122_cse | or_188_cse;
  assign or_dcpl_50 = (~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4);
  assign or_dcpl_53 = (~ or_185_cse) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4);
  assign and_dcpl_123 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]));
  assign and_dcpl_124 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]));
  assign and_dcpl_125 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]));
  assign and_dcpl_126 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]));
  assign and_dcpl_127 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]));
  assign and_dcpl_128 = (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]) & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]));
  assign and_dcpl_129 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign and_dcpl_130 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign and_dcpl_133 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_137 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign and_dcpl_154 = and_dcpl_133 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]);
  assign and_dcpl_155 = and_dcpl_133 & and_dcpl_123;
  assign and_dcpl_156 = and_dcpl_133 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]);
  assign and_dcpl_157 = and_dcpl_133 & and_dcpl_128;
  assign and_dcpl_158 = and_dcpl_133 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]);
  assign and_dcpl_159 = and_dcpl_133 & and_dcpl_127;
  assign and_dcpl_160 = and_dcpl_133 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]);
  assign and_dcpl_161 = and_dcpl_133 & and_dcpl_125;
  assign and_dcpl_162 = and_dcpl_133 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]);
  assign and_dcpl_163 = and_dcpl_133 & and_dcpl_126;
  assign and_dcpl_164 = and_dcpl_133 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]);
  assign and_dcpl_165 = and_dcpl_133 & and_dcpl_124;
  assign and_dcpl_166 = and_dcpl_133 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]);
  assign and_dcpl_167 = and_dcpl_133 & and_dcpl_129;
  assign and_dcpl_168 = and_dcpl_133 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]);
  assign and_dcpl_169 = and_dcpl_133 & and_dcpl_130;
  assign and_dcpl_172 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign and_dcpl_176 = (state_2_1_sva==2'b01) & (~ state_0_sva) & and_626_cse;
  assign mux_10_nl = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      state_2_1_sva[1]);
  assign and_753_nl = (state_2_1_sva[1]) & PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  assign mux_11_nl = MUX_s_1_2_2(mux_10_nl, and_753_nl, state_2_1_sva[0]);
  assign mux_12_nl = MUX_s_1_2_2(mux_11_nl, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      state_0_sva);
  assign and_dcpl_179 = mux_12_nl & (~(PECore_RunFSM_switch_lp_nor_tmp_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign and_dcpl_180 = rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign or_dcpl_121 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]!=2'b01);
  assign or_dcpl_126 = ~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_129 = or_dcpl_121 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign and_dcpl_183 = reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign and_dcpl_186 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01);
  assign and_dcpl_187 = and_dcpl_186 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]))
      & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign and_dcpl_188 = and_dcpl_187 & and_dcpl_183 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_189 = reg_rva_in_PopNB_mioi_iswt0_cse & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_191 = and_dcpl_187 & and_dcpl_189 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_195 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7;
  assign or_tmp_35 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      | rva_in_reg_rw_sva_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1
      | rva_in_reg_rw_sva_st_1_4;
  assign and_dcpl_226 = and_dcpl_180 & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_230 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9
      & (~ rva_in_reg_rw_sva_st_1_9);
  assign and_dcpl_231 = and_dcpl_230 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign and_dcpl_241 = ~(input_read_req_valid_lpi_1_dfm_1_9 | rva_in_reg_rw_sva_9);
  assign and_dcpl_253 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1;
  assign and_dcpl_258 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & while_stage_0_6;
  assign not_tmp_139 = ~(rva_in_reg_rw_sva_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1
      | rva_in_reg_rw_sva_st_1_4);
  assign nand_29_nl = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign or_203_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])
      | (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_45_nl = MUX_s_1_2_2(nand_29_nl, or_203_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign or_202_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]!=2'b00)
      | (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign mux_tmp_46 = MUX_s_1_2_2(mux_45_nl, or_202_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign and_dcpl_274 = PECore_RunFSM_switch_lp_equal_tmp_1_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_282 = and_dcpl_186 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]))
      & and_dcpl_180;
  assign and_dcpl_284 = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_5);
  assign and_dcpl_312 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
      & (~ rva_in_reg_rw_sva_st_1_8);
  assign and_dcpl_313 = and_dcpl_312 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6);
  assign and_dcpl_320 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      & while_stage_0_8;
  assign and_dcpl_321 = PECore_RunMac_PECore_RunMac_if_and_svs_st_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign and_759_nl = (Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3_1 |
      Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp)
      & PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign mux_tmp_51 = MUX_s_1_2_2(and_759_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3_1);
  assign or_tmp_59 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ mux_tmp_51);
  assign and_dcpl_325 = ~(rva_in_reg_rw_sva_8 | input_read_req_valid_lpi_1_dfm_1_8);
  assign and_dcpl_343 = (~ rva_in_reg_rw_sva_st_1_7) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  assign and_dcpl_344 = and_dcpl_343 & while_stage_0_9;
  assign and_dcpl_347 = while_stage_0_9 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5)
      & (~ input_read_req_valid_lpi_1_dfm_1_7);
  assign and_dcpl_348 = PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 & (~ rva_in_reg_rw_sva_7);
  assign or_dcpl_177 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:2]!=2'b00);
  assign or_dcpl_178 = or_dcpl_177 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]);
  assign or_dcpl_179 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]!=2'b00);
  assign or_dcpl_180 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]);
  assign or_dcpl_181 = or_dcpl_180 | or_dcpl_179;
  assign or_dcpl_182 = or_dcpl_181 | or_dcpl_178;
  assign or_dcpl_185 = or_dcpl_129 | or_dcpl_126 | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]);
  assign or_dcpl_187 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]!=2'b01);
  assign or_dcpl_188 = or_dcpl_180 | or_dcpl_187;
  assign or_dcpl_189 = or_dcpl_188 | or_dcpl_178;
  assign or_dcpl_191 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]!=2'b10);
  assign or_dcpl_192 = or_dcpl_180 | or_dcpl_191;
  assign or_dcpl_193 = or_dcpl_192 | or_dcpl_178;
  assign or_dcpl_195 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]==2'b11));
  assign or_dcpl_196 = or_dcpl_180 | or_dcpl_195;
  assign or_dcpl_197 = or_dcpl_196 | or_dcpl_178;
  assign or_dcpl_199 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:2]!=2'b01);
  assign or_dcpl_200 = or_dcpl_199 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]);
  assign or_dcpl_201 = or_dcpl_181 | or_dcpl_200;
  assign or_dcpl_203 = or_dcpl_188 | or_dcpl_200;
  assign or_dcpl_205 = or_dcpl_192 | or_dcpl_200;
  assign or_dcpl_207 = or_dcpl_196 | or_dcpl_200;
  assign or_dcpl_209 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:2]!=2'b10);
  assign or_dcpl_210 = or_dcpl_209 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]);
  assign or_dcpl_211 = or_dcpl_181 | or_dcpl_210;
  assign or_dcpl_213 = or_dcpl_188 | or_dcpl_210;
  assign or_dcpl_215 = or_dcpl_192 | or_dcpl_210;
  assign or_dcpl_217 = or_dcpl_196 | or_dcpl_210;
  assign or_dcpl_219 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:2]==2'b11));
  assign or_dcpl_220 = or_dcpl_219 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]);
  assign or_dcpl_221 = or_dcpl_181 | or_dcpl_220;
  assign or_dcpl_223 = or_dcpl_188 | or_dcpl_220;
  assign or_dcpl_225 = or_dcpl_192 | or_dcpl_220;
  assign or_dcpl_227 = or_dcpl_196 | or_dcpl_220;
  assign or_dcpl_229 = or_dcpl_177 | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]));
  assign or_dcpl_230 = or_dcpl_181 | or_dcpl_229;
  assign or_dcpl_232 = or_dcpl_188 | or_dcpl_229;
  assign or_dcpl_234 = or_dcpl_192 | or_dcpl_229;
  assign or_dcpl_236 = or_dcpl_196 | or_dcpl_229;
  assign or_dcpl_238 = or_dcpl_199 | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]));
  assign or_dcpl_239 = or_dcpl_181 | or_dcpl_238;
  assign or_dcpl_241 = or_dcpl_188 | or_dcpl_238;
  assign or_dcpl_243 = or_dcpl_192 | or_dcpl_238;
  assign or_dcpl_245 = or_dcpl_196 | or_dcpl_238;
  assign or_dcpl_247 = or_dcpl_209 | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]));
  assign or_dcpl_248 = or_dcpl_181 | or_dcpl_247;
  assign or_dcpl_250 = or_dcpl_188 | or_dcpl_247;
  assign or_dcpl_252 = or_dcpl_192 | or_dcpl_247;
  assign or_dcpl_254 = or_dcpl_196 | or_dcpl_247;
  assign or_dcpl_256 = or_dcpl_219 | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]));
  assign or_dcpl_257 = or_dcpl_181 | or_dcpl_256;
  assign or_dcpl_259 = or_dcpl_188 | or_dcpl_256;
  assign or_dcpl_261 = or_dcpl_192 | or_dcpl_256;
  assign or_dcpl_263 = or_dcpl_196 | or_dcpl_256;
  assign or_dcpl_265 = (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]);
  assign or_dcpl_266 = or_dcpl_265 | or_dcpl_179;
  assign or_dcpl_267 = or_dcpl_266 | or_dcpl_178;
  assign or_dcpl_269 = or_dcpl_265 | or_dcpl_187;
  assign or_dcpl_270 = or_dcpl_269 | or_dcpl_178;
  assign or_dcpl_272 = or_dcpl_265 | or_dcpl_191;
  assign or_dcpl_273 = or_dcpl_272 | or_dcpl_178;
  assign or_dcpl_275 = or_dcpl_265 | or_dcpl_195;
  assign or_dcpl_276 = or_dcpl_275 | or_dcpl_178;
  assign or_dcpl_278 = or_dcpl_266 | or_dcpl_200;
  assign or_dcpl_280 = or_dcpl_269 | or_dcpl_200;
  assign or_dcpl_282 = or_dcpl_272 | or_dcpl_200;
  assign or_dcpl_284 = or_dcpl_275 | or_dcpl_200;
  assign or_dcpl_286 = or_dcpl_266 | or_dcpl_210;
  assign or_dcpl_288 = or_dcpl_269 | or_dcpl_210;
  assign or_dcpl_290 = or_dcpl_272 | or_dcpl_210;
  assign or_dcpl_292 = or_dcpl_275 | or_dcpl_210;
  assign or_dcpl_294 = or_dcpl_266 | or_dcpl_220;
  assign or_dcpl_296 = or_dcpl_269 | or_dcpl_220;
  assign or_dcpl_298 = or_dcpl_272 | or_dcpl_220;
  assign or_dcpl_300 = or_dcpl_275 | or_dcpl_220;
  assign or_dcpl_302 = or_dcpl_266 | or_dcpl_229;
  assign or_dcpl_304 = or_dcpl_269 | or_dcpl_229;
  assign or_dcpl_306 = or_dcpl_272 | or_dcpl_229;
  assign or_dcpl_308 = or_dcpl_275 | or_dcpl_229;
  assign or_dcpl_310 = or_dcpl_266 | or_dcpl_238;
  assign or_dcpl_312 = or_dcpl_269 | or_dcpl_238;
  assign or_dcpl_314 = or_dcpl_272 | or_dcpl_238;
  assign or_dcpl_316 = or_dcpl_275 | or_dcpl_238;
  assign or_dcpl_318 = or_dcpl_266 | or_dcpl_247;
  assign or_dcpl_320 = or_dcpl_269 | or_dcpl_247;
  assign or_dcpl_322 = or_dcpl_272 | or_dcpl_247;
  assign or_dcpl_324 = or_dcpl_275 | or_dcpl_247;
  assign or_dcpl_326 = or_dcpl_266 | or_dcpl_256;
  assign or_dcpl_328 = or_dcpl_269 | or_dcpl_256;
  assign or_dcpl_330 = or_dcpl_272 | or_dcpl_256;
  assign or_dcpl_332 = or_dcpl_275 | or_dcpl_256;
  assign or_dcpl_336 = or_dcpl_129 | or_dcpl_126 | (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])));
  assign or_dcpl_401 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]));
  assign or_dcpl_402 = or_dcpl_401 | or_dcpl_179;
  assign or_dcpl_403 = or_dcpl_402 | or_dcpl_178;
  assign or_dcpl_405 = or_dcpl_401 | or_dcpl_187;
  assign or_dcpl_406 = or_dcpl_405 | or_dcpl_178;
  assign or_dcpl_408 = or_dcpl_401 | or_dcpl_191;
  assign or_dcpl_409 = or_dcpl_408 | or_dcpl_178;
  assign or_dcpl_411 = or_dcpl_401 | or_dcpl_195;
  assign or_dcpl_412 = or_dcpl_411 | or_dcpl_178;
  assign or_dcpl_414 = or_dcpl_402 | or_dcpl_200;
  assign or_dcpl_416 = or_dcpl_405 | or_dcpl_200;
  assign or_dcpl_418 = or_dcpl_408 | or_dcpl_200;
  assign or_dcpl_420 = or_dcpl_411 | or_dcpl_200;
  assign or_dcpl_422 = or_dcpl_402 | or_dcpl_210;
  assign or_dcpl_424 = or_dcpl_405 | or_dcpl_210;
  assign or_dcpl_426 = or_dcpl_408 | or_dcpl_210;
  assign or_dcpl_428 = or_dcpl_411 | or_dcpl_210;
  assign or_dcpl_430 = or_dcpl_402 | or_dcpl_220;
  assign or_dcpl_432 = or_dcpl_405 | or_dcpl_220;
  assign or_dcpl_434 = or_dcpl_408 | or_dcpl_220;
  assign or_dcpl_436 = or_dcpl_411 | or_dcpl_220;
  assign or_dcpl_438 = or_dcpl_402 | or_dcpl_229;
  assign or_dcpl_440 = or_dcpl_405 | or_dcpl_229;
  assign or_dcpl_442 = or_dcpl_408 | or_dcpl_229;
  assign or_dcpl_444 = or_dcpl_411 | or_dcpl_229;
  assign or_dcpl_446 = or_dcpl_402 | or_dcpl_238;
  assign or_dcpl_448 = or_dcpl_405 | or_dcpl_238;
  assign or_dcpl_450 = or_dcpl_408 | or_dcpl_238;
  assign or_dcpl_452 = or_dcpl_411 | or_dcpl_238;
  assign or_dcpl_454 = or_dcpl_402 | or_dcpl_247;
  assign or_dcpl_456 = or_dcpl_405 | or_dcpl_247;
  assign or_dcpl_458 = or_dcpl_408 | or_dcpl_247;
  assign or_dcpl_460 = or_dcpl_411 | or_dcpl_247;
  assign or_dcpl_462 = or_dcpl_402 | or_dcpl_256;
  assign or_dcpl_464 = or_dcpl_405 | or_dcpl_256;
  assign or_dcpl_466 = or_dcpl_408 | or_dcpl_256;
  assign or_dcpl_468 = or_dcpl_411 | or_dcpl_256;
  assign or_dcpl_470 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]));
  assign or_dcpl_471 = or_dcpl_470 | or_dcpl_179;
  assign or_dcpl_472 = or_dcpl_471 | or_dcpl_178;
  assign or_dcpl_474 = or_dcpl_470 | or_dcpl_187;
  assign or_dcpl_475 = or_dcpl_474 | or_dcpl_178;
  assign or_dcpl_477 = or_dcpl_470 | or_dcpl_191;
  assign or_dcpl_478 = or_dcpl_477 | or_dcpl_178;
  assign or_dcpl_480 = or_dcpl_470 | or_dcpl_195;
  assign or_dcpl_481 = or_dcpl_480 | or_dcpl_178;
  assign or_dcpl_483 = or_dcpl_471 | or_dcpl_200;
  assign or_dcpl_485 = or_dcpl_474 | or_dcpl_200;
  assign or_dcpl_487 = or_dcpl_477 | or_dcpl_200;
  assign or_dcpl_489 = or_dcpl_480 | or_dcpl_200;
  assign or_dcpl_491 = or_dcpl_471 | or_dcpl_210;
  assign or_dcpl_493 = or_dcpl_474 | or_dcpl_210;
  assign or_dcpl_495 = or_dcpl_477 | or_dcpl_210;
  assign or_dcpl_497 = or_dcpl_480 | or_dcpl_210;
  assign or_dcpl_499 = or_dcpl_471 | or_dcpl_220;
  assign or_dcpl_501 = or_dcpl_474 | or_dcpl_220;
  assign or_dcpl_503 = or_dcpl_477 | or_dcpl_220;
  assign or_dcpl_505 = or_dcpl_480 | or_dcpl_220;
  assign or_dcpl_507 = or_dcpl_471 | or_dcpl_229;
  assign or_dcpl_509 = or_dcpl_474 | or_dcpl_229;
  assign or_dcpl_511 = or_dcpl_477 | or_dcpl_229;
  assign or_dcpl_513 = or_dcpl_480 | or_dcpl_229;
  assign or_dcpl_515 = or_dcpl_471 | or_dcpl_238;
  assign or_dcpl_517 = or_dcpl_474 | or_dcpl_238;
  assign or_dcpl_519 = or_dcpl_477 | or_dcpl_238;
  assign or_dcpl_521 = or_dcpl_480 | or_dcpl_238;
  assign or_dcpl_523 = or_dcpl_471 | or_dcpl_247;
  assign or_dcpl_525 = or_dcpl_474 | or_dcpl_247;
  assign or_dcpl_527 = or_dcpl_477 | or_dcpl_247;
  assign or_dcpl_529 = or_dcpl_480 | or_dcpl_247;
  assign or_dcpl_531 = or_dcpl_471 | or_dcpl_256;
  assign or_dcpl_533 = or_dcpl_474 | or_dcpl_256;
  assign or_dcpl_535 = or_dcpl_477 | or_dcpl_256;
  assign or_dcpl_537 = or_dcpl_480 | or_dcpl_256;
  assign and_dcpl_367 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & while_stage_0_8;
  assign and_dcpl_371 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & (~ rva_in_reg_rw_sva_st_1_6);
  assign and_dcpl_372 = and_dcpl_371 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4);
  assign and_dcpl_380 = ~(rva_in_reg_rw_sva_6 | input_read_req_valid_lpi_1_dfm_1_6);
  assign and_dcpl_395 = while_stage_0_7 & (~ rva_in_reg_rw_sva_st_1_5);
  assign and_dcpl_408 = while_and_21_cse & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_dcpl_423 = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)
      & while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign and_dcpl_444 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1
      | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_363_itm_1);
  assign or_tmp_68 = input_read_req_valid_lpi_1_dfm_1_3 | rva_in_reg_rw_sva_3 | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_363_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign and_dcpl_457 = and_dcpl_444 & (~ rva_in_reg_rw_sva_3);
  assign or_dcpl_606 = (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp)
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_tmp;
  assign and_dcpl_468 = or_dcpl_606 & (~(reg_rva_in_reg_rw_sva_2_cse | input_read_req_valid_lpi_1_dfm_1_2));
  assign and_dcpl_488 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | input_read_req_valid_lpi_1_dfm_1_1);
  assign and_dcpl_489 = and_dcpl_488 & and_dcpl_172;
  assign mux_tmp_69 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1!=4'b0100));
  assign and_dcpl_495 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1);
  assign nand_35_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) & PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp);
  assign and_dcpl_530 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_7 & while_stage_0_9;
  assign and_dcpl_532 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_6 & while_stage_0_8;
  assign or_tmp_75 = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9) | (~ while_stage_0_11)
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_9 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9;
  assign or_tmp_76 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_10
      | (~ while_stage_0_12);
  assign or_tmp_78 = PECore_RunMac_PECore_RunMac_if_and_svs_st_9 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9;
  assign and_dcpl_544 = and_dcpl_76 & (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]);
  assign or_698_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1;
  assign mux_74_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      or_698_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_tmp_2 = while_stage_0_6 & mux_74_nl;
  assign and_dcpl_546 = and_dcpl_76 & (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign or_702_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_1;
  assign mux_77_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      or_702_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_tmp_3 = while_stage_0_6 & mux_77_nl;
  assign or_708_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]);
  assign mux_83_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_708_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_4 = while_stage_0_5 & mux_83_nl;
  assign or_713_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_380_itm_1
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]);
  assign mux_86_nl = MUX_s_1_2_2(or_50_cse, or_713_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_5 = while_stage_0_5 & mux_86_nl;
  assign or_721_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]);
  assign mux_89_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_721_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_6 = while_stage_0_5 & mux_89_nl;
  assign or_724_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_3 | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]);
  assign mux_92_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_724_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_7 = while_stage_0_5 & mux_92_nl;
  assign or_732_nl = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp
      | (or_dcpl_32 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign mux_95_nl = MUX_s_1_2_2(or_732_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse);
  assign or_tmp_111 = Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp
      | mux_95_nl;
  assign or_728_nl = PECore_UpdateFSM_switch_lp_equal_tmp_2_3 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  assign mux_96_nl = MUX_s_1_2_2(or_tmp_111, or_728_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_8 = while_stage_0_5 & mux_96_nl;
  assign or_738_nl = PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 | PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign mux_99_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_738_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_tmp_9 = while_stage_0_5 & mux_99_nl;
  assign and_dcpl_567 = fsm_output & (~ weight_mem_run_3_for_land_5_lpi_1_dfm_3);
  assign and_dcpl_568 = fsm_output & (~ weight_mem_run_3_for_land_3_lpi_1_dfm_3);
  assign or_dcpl_633 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7);
  assign and_dcpl_584 = (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) |
      (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]))) & nor_279_cse;
  assign and_dcpl_588 = nor_276_cse & (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]))) & and_dcpl_584;
  assign and_dcpl_590 = (~(while_stage_0_4 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
      & while_stage_0_5;
  assign or_dcpl_636 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ while_stage_0_5);
  assign or_dcpl_637 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ while_stage_0_3);
  assign or_dcpl_648 = nand_83_cse | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_649 = or_dcpl_121 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]);
  assign and_dcpl_621 = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) |
      (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]));
  assign and_dcpl_635 = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]) |
      (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]));
  assign or_dcpl_700 = (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | nand_35_cse;
  assign and_dcpl_657 = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2:1]==2'b10);
  assign and_dcpl_664 = ~(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign and_dcpl_674 = weight_mem_run_3_for_land_7_lpi_1_dfm_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_dcpl_675 = ~(weight_mem_run_3_for_land_7_lpi_1_dfm_2 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_dcpl_706 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      | rva_in_reg_rw_sva_6 | (~ while_stage_0_8);
  assign and_777_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]) & while_mux_1471_tmp;
  assign and_778_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) & while_mux_1473_tmp;
  assign or_tmp_131 = and_777_cse | and_778_cse;
  assign and_779_cse = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1;
  assign and_780_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  assign or_tmp_133 = and_779_cse | and_780_cse;
  assign mux_125_nl = MUX_s_1_2_2(or_tmp_133, or_tmp_131, while_stage_0_5);
  assign or_843_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva | or_tmp_133;
  assign or_841_nl = while_mux_1472_tmp | or_tmp_131;
  assign mux_124_nl = MUX_s_1_2_2(or_843_nl, or_841_nl, while_stage_0_5);
  assign mux_tmp_126 = MUX_s_1_2_2(mux_125_nl, mux_124_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign nor_tmp_45 = while_mux_1476_tmp & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign and_782_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) & while_mux_1477_tmp;
  assign or_tmp_135 = and_782_cse | nor_tmp_45;
  assign and_783_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) & while_mux_1474_tmp;
  assign or_tmp_136 = and_783_cse | or_tmp_135;
  assign and_784_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) & while_mux_1475_tmp;
  assign or_tmp_137 = and_784_cse | or_tmp_136;
  assign or_tmp_139 = and_777_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])
      & while_mux_1473_tmp)) & or_tmp_137));
  assign nor_tmp_51 = weight_mem_read_arbxbar_arbiters_next_7_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign and_788_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  assign or_tmp_141 = and_788_cse | nor_tmp_51;
  assign and_789_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  assign or_tmp_142 = and_789_cse | or_tmp_141;
  assign and_790_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  assign or_tmp_143 = and_790_cse | or_tmp_142;
  assign or_tmp_145 = and_779_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])
      & weight_mem_read_arbxbar_arbiters_next_7_5_sva)) & or_tmp_143));
  assign mux_128_nl = MUX_s_1_2_2(or_tmp_145, or_tmp_139, while_stage_0_5);
  assign or_855_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva | or_tmp_145;
  assign or_849_nl = while_mux_1472_tmp | or_tmp_139;
  assign mux_127_nl = MUX_s_1_2_2(or_855_nl, or_849_nl, while_stage_0_5);
  assign mux_129_itm = MUX_s_1_2_2(mux_128_nl, mux_127_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign or_tmp_149 = and_782_cse | nor_tmp_45 | and_784_cse | and_783_cse;
  assign or_tmp_150 = and_778_cse | or_tmp_149;
  assign or_tmp_151 = and_777_cse | or_tmp_150;
  assign or_tmp_155 = and_788_cse | nor_tmp_51 | and_790_cse | and_789_cse;
  assign or_tmp_156 = and_780_cse | or_tmp_155;
  assign or_tmp_157 = and_779_cse | or_tmp_156;
  assign or_873_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])) | weight_mem_read_arbxbar_arbiters_next_7_5_sva
      | or_tmp_155;
  assign or_871_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | or_tmp_156;
  assign mux_133_nl = MUX_s_1_2_2(or_873_nl, or_871_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign mux_134_nl = MUX_s_1_2_2(mux_133_nl, or_tmp_157, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign or_870_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])) | while_mux_1473_tmp
      | or_tmp_149;
  assign or_868_nl = while_mux_1471_tmp | or_tmp_150;
  assign mux_131_nl = MUX_s_1_2_2(or_870_nl, or_868_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign mux_132_nl = MUX_s_1_2_2(mux_131_nl, or_tmp_151, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign mux_135_nl = MUX_s_1_2_2(mux_134_nl, mux_132_nl, while_stage_0_5);
  assign or_867_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva | or_tmp_157;
  assign or_861_nl = while_mux_1472_tmp | or_tmp_151;
  assign mux_130_nl = MUX_s_1_2_2(or_867_nl, or_861_nl, while_stage_0_5);
  assign mux_136_itm = MUX_s_1_2_2(mux_135_nl, mux_130_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign nor_384_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_2_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])));
  assign nor_385_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_1_sva | nor_tmp_51);
  assign mux_140_nl = MUX_s_1_2_2(nor_384_nl, nor_385_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign nor_386_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_4_sva | or_tmp_141);
  assign mux_141_nl = MUX_s_1_2_2(mux_140_nl, nor_386_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign nor_387_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_3_sva | or_tmp_142);
  assign mux_142_nl = MUX_s_1_2_2(mux_141_nl, nor_387_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nor_388_nl = ~(while_mux_1476_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])));
  assign nor_389_nl = ~(while_mux_1477_tmp | nor_tmp_45);
  assign mux_137_nl = MUX_s_1_2_2(nor_388_nl, nor_389_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign nor_390_nl = ~(while_mux_1474_tmp | or_tmp_135);
  assign mux_138_nl = MUX_s_1_2_2(mux_137_nl, nor_390_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign nor_391_nl = ~(while_mux_1475_tmp | or_tmp_136);
  assign mux_139_nl = MUX_s_1_2_2(mux_138_nl, nor_391_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign mux_143_nl = MUX_s_1_2_2(mux_142_nl, mux_139_nl, while_stage_0_5);
  assign and_dcpl_680 = mux_143_nl & and_dcpl_584;
  assign or_tmp_174 = and_777_cse | and_778_cse | or_tmp_137;
  assign or_tmp_177 = and_779_cse | and_780_cse | or_tmp_143;
  assign and_810_cse = while_mux_1464_tmp & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_tmp_179 = ((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & while_mux_1466_tmp)
      | and_810_cse;
  assign or_tmp_181 = ((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_5_sva)
      | (Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]));
  assign mux_148_nl = MUX_s_1_2_2(or_tmp_181, or_tmp_179, while_stage_0_5);
  assign or_891_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | or_tmp_181;
  assign or_889_nl = while_mux_1465_tmp | or_tmp_179;
  assign mux_147_nl = MUX_s_1_2_2(or_891_nl, or_889_nl, while_stage_0_5);
  assign mux_tmp_149 = MUX_s_1_2_2(mux_148_nl, mux_147_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign and_814_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & while_mux_1469_tmp;
  assign and_815_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) & while_mux_1467_tmp;
  assign and_816_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & while_mux_1468_tmp;
  assign nand_6_nl = ~(while_mux_1470_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      & (~ or_tmp_179));
  assign mux_150_nl = MUX_s_1_2_2(nand_6_nl, or_tmp_179, and_814_cse);
  assign mux_151_nl = MUX_s_1_2_2(mux_150_nl, or_tmp_179, and_815_cse);
  assign mux_tmp_152 = MUX_s_1_2_2(mux_151_nl, or_tmp_179, and_816_cse);
  assign and_818_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  assign and_819_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  assign and_820_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  assign nand_7_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      & (~ or_tmp_181));
  assign mux_153_nl = MUX_s_1_2_2(nand_7_nl, or_tmp_181, and_818_cse);
  assign mux_154_nl = MUX_s_1_2_2(mux_153_nl, or_tmp_181, and_819_cse);
  assign mux_tmp_155 = MUX_s_1_2_2(mux_154_nl, or_tmp_181, and_820_cse);
  assign mux_157_nl = MUX_s_1_2_2(mux_tmp_155, mux_tmp_152, while_stage_0_5);
  assign or_893_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | mux_tmp_155;
  assign or_892_nl = while_mux_1465_tmp | mux_tmp_152;
  assign mux_156_nl = MUX_s_1_2_2(or_893_nl, or_892_nl, while_stage_0_5);
  assign mux_158_itm = MUX_s_1_2_2(mux_157_nl, mux_156_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign nor_tmp_83 = while_mux_1465_tmp & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign or_tmp_186 = and_810_cse | nor_tmp_83;
  assign or_898_nl = while_mux_1465_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign or_897_nl = while_mux_1464_tmp | nor_tmp_83;
  assign mux_159_nl = MUX_s_1_2_2(or_898_nl, or_897_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_160_nl = MUX_s_1_2_2(mux_159_nl, or_tmp_186, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_896_nl = while_mux_1466_tmp | or_tmp_186;
  assign mux_161_nl = MUX_s_1_2_2(mux_160_nl, or_896_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_191 = and_814_cse | and_815_cse | mux_161_nl;
  assign and_825_cse = weight_mem_read_arbxbar_arbiters_next_6_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign or_tmp_194 = and_825_cse | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  assign mux_tmp_162 = MUX_s_1_2_2(and_825_cse, or_tmp_194, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_905_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign mux_163_nl = MUX_s_1_2_2(or_905_nl, or_tmp_194, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_164_nl = MUX_s_1_2_2(mux_163_nl, mux_tmp_162, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_904_nl = weight_mem_read_arbxbar_arbiters_next_6_5_sva | mux_tmp_162;
  assign mux_165_nl = MUX_s_1_2_2(mux_164_nl, or_904_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_198 = and_818_cse | and_819_cse | mux_165_nl;
  assign mux_170_nl = MUX_s_1_2_2(or_tmp_198, or_tmp_191, while_stage_0_5);
  assign or_912_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | or_tmp_198;
  assign or_911_nl = while_mux_1468_tmp | or_tmp_191;
  assign mux_169_nl = MUX_s_1_2_2(or_912_nl, or_911_nl, while_stage_0_5);
  assign mux_171_nl = MUX_s_1_2_2(mux_170_nl, mux_169_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign or_910_nl = weight_mem_read_arbxbar_arbiters_next_6_1_sva | or_tmp_198;
  assign or_909_nl = while_mux_1470_tmp | or_tmp_191;
  assign mux_167_nl = MUX_s_1_2_2(or_910_nl, or_909_nl, while_stage_0_5);
  assign or_908_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | or_tmp_198;
  assign or_901_nl = while_mux_1468_tmp | while_mux_1470_tmp | or_tmp_191;
  assign mux_166_nl = MUX_s_1_2_2(or_908_nl, or_901_nl, while_stage_0_5);
  assign mux_168_nl = MUX_s_1_2_2(mux_167_nl, mux_166_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_172_itm = MUX_s_1_2_2(mux_171_nl, mux_168_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign nor_tmp_90 = while_mux_1470_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_tmp_204 = and_814_cse | nor_tmp_90;
  assign nor_tmp_93 = weight_mem_read_arbxbar_arbiters_next_6_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_tmp_210 = and_818_cse | nor_tmp_93;
  assign nor_392_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_1_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])));
  assign nor_393_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_2_sva | nor_tmp_93);
  assign mux_176_nl = MUX_s_1_2_2(nor_392_nl, nor_393_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign nor_394_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_4_sva | or_tmp_210);
  assign mux_177_nl = MUX_s_1_2_2(mux_176_nl, nor_394_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign nor_395_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_3_sva | and_819_cse
      | or_tmp_210);
  assign mux_178_nl = MUX_s_1_2_2(mux_177_nl, nor_395_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nor_396_nl = ~(while_mux_1470_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])));
  assign nor_397_nl = ~(while_mux_1469_tmp | nor_tmp_90);
  assign mux_173_nl = MUX_s_1_2_2(nor_396_nl, nor_397_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign nor_398_nl = ~(while_mux_1467_tmp | or_tmp_204);
  assign mux_174_nl = MUX_s_1_2_2(mux_173_nl, nor_398_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign nor_399_nl = ~(while_mux_1468_tmp | and_815_cse | or_tmp_204);
  assign mux_175_nl = MUX_s_1_2_2(mux_174_nl, nor_399_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_179_nl = MUX_s_1_2_2(mux_178_nl, mux_175_nl, while_stage_0_5);
  assign and_dcpl_683 = mux_179_nl & nor_280_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6])));
  assign or_tmp_219 = and_816_cse | and_815_cse | and_814_cse | nor_tmp_90 | or_tmp_179;
  assign or_tmp_224 = and_820_cse | and_819_cse | and_818_cse | nor_tmp_93 | or_tmp_181;
  assign while_mux_1482_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_183_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1,
      while_mux_1482_nl, while_stage_0_5);
  assign or_dcpl_710 = (mux_183_nl & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]))
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  assign and_dcpl_685 = ~(weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp);
  assign Arbiter_8U_Roundrobin_pick_1_mux_595_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1463_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_595_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_843_cse = while_mux_1463_nl & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign or_tmp_226 = and_843_cse | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp;
  assign and_844_cse = weight_mem_read_arbxbar_arbiters_next_5_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign or_tmp_228 = and_844_cse | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp;
  assign mux_185_nl = MUX_s_1_2_2(or_tmp_228, or_tmp_226, while_stage_0_5);
  assign nor_402_nl = ~(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1
      | (~ or_tmp_228));
  assign nor_403_nl = ~(while_mux_1457_cse_1 | (~ or_tmp_226));
  assign mux_184_nl = MUX_s_1_2_2(nor_402_nl, nor_403_nl, while_stage_0_5);
  assign mux_186_nl = MUX_s_1_2_2(mux_185_nl, mux_184_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign and_dcpl_686 = mux_186_nl & and_dcpl_685;
  assign and_dcpl_687 = ~(weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp);
  assign and_dcpl_688 = and_dcpl_685 & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp);
  assign and_dcpl_689 = and_dcpl_688 & and_dcpl_687;
  assign or_943_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1
      | and_844_cse;
  assign or_942_nl = while_mux_1457_cse_1 | and_843_cse;
  assign mux_tmp_187 = MUX_s_1_2_2(or_943_nl, or_942_nl, while_stage_0_5);
  assign mux_tmp_188 = MUX_s_1_2_2(and_844_cse, and_843_cse, while_stage_0_5);
  assign mux_tmp_189 = MUX_s_1_2_2(mux_tmp_188, mux_tmp_187, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign nand_8_nl = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) & (~
      mux_tmp_188));
  assign mux_190_nl = MUX_s_1_2_2(nand_8_nl, mux_tmp_187, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign or_941_nl = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign mux_191_nl = MUX_s_1_2_2(mux_190_nl, mux_tmp_189, or_941_nl);
  assign and_dcpl_690 = (~ mux_191_nl) & and_dcpl_689;
  assign and_dcpl_696 = (~ mux_tmp_188) & and_dcpl_688 & and_dcpl_687 & (~ (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]))
      & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5])));
  assign nor_tmp_107 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]) & while_mux_1450_tmp;
  assign nor_tmp_109 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1;
  assign or_944_cse = and_999_cse | nor_tmp_107;
  assign or_945_cse = and_997_cse | nor_tmp_109;
  assign mux_192_cse = MUX_s_1_2_2(or_945_cse, or_944_cse, while_stage_0_5);
  assign or_dcpl_711 = mux_192_cse | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign nand_tmp_9 = ~(while_mux_1456_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      & (~ or_944_cse));
  assign nand_tmp_10 = ~(weight_mem_read_arbxbar_arbiters_next_4_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      & (~ or_945_cse));
  assign mux_197_nl = MUX_s_1_2_2(nand_tmp_10, nand_tmp_9, while_stage_0_5);
  assign mux_195_nl = MUX_s_1_2_2(nand_tmp_10, or_945_cse, weight_mem_read_arbxbar_arbiters_next_4_3_sva);
  assign mux_194_nl = MUX_s_1_2_2(nand_tmp_9, or_944_cse, while_mux_1454_tmp);
  assign mux_196_nl = MUX_s_1_2_2(mux_195_nl, mux_194_nl, while_stage_0_5);
  assign mux_198_nl = MUX_s_1_2_2(mux_197_nl, mux_196_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign or_947_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  assign mux_199_nl = MUX_s_1_2_2(mux_198_nl, mux_192_cse, or_947_nl);
  assign and_dcpl_698 = ~(mux_199_nl | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp);
  assign and_dcpl_700 = ~(weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp);
  assign and_857_cse = while_mux_1456_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign or_tmp_238 = and_857_cse | nor_tmp_107;
  assign and_858_cse = weight_mem_read_arbxbar_arbiters_next_4_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign or_tmp_242 = and_858_cse | nor_tmp_109;
  assign mux_202_nl = MUX_s_1_2_2(nor_284_cse, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1,
      weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign or_956_nl = and_858_cse | mux_202_nl;
  assign or_955_nl = weight_mem_read_arbxbar_arbiters_next_4_6_sva | or_tmp_242;
  assign mux_203_nl = MUX_s_1_2_2(or_956_nl, or_955_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign nor_410_nl = ~(and_996_cse | mux_203_nl);
  assign mux_200_nl = MUX_s_1_2_2(nor_284_cse, while_mux_1450_tmp, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign or_952_nl = and_857_cse | mux_200_nl;
  assign or_951_nl = while_mux_1451_tmp | or_tmp_238;
  assign mux_201_nl = MUX_s_1_2_2(or_952_nl, or_951_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign nor_411_nl = ~(and_998_cse | mux_201_nl);
  assign mux_204_nl = MUX_s_1_2_2(nor_410_nl, nor_411_nl, while_stage_0_5);
  assign and_dcpl_701 = mux_204_nl & and_dcpl_700;
  assign nor_412_nl = ~(and_996_cse | and_858_cse);
  assign nor_413_nl = ~(and_998_cse | and_857_cse);
  assign mux_205_nl = MUX_s_1_2_2(nor_412_nl, nor_413_nl, while_stage_0_5);
  assign and_dcpl_707 = mux_205_nl & nor_284_cse & (~(weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4])
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp));
  assign mux_207_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_5_sva,
      while_mux_1445_tmp, while_stage_0_5);
  assign or_dcpl_713 = (mux_207_nl & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]))
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_mux_610_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1446_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_610_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_867_cse = while_mux_1446_nl & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign or_tmp_253 = and_867_cse | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  assign nor_tmp_135 = ~(Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1));
  assign nor_tmp_136 = Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign or_975_nl = nor_tmp_136 | or_tmp_253;
  assign nand_12_nl = ~(nor_tmp_135 & (~ or_tmp_253));
  assign mux_210_nl = MUX_s_1_2_2(or_975_nl, nand_12_nl, weight_mem_read_arbxbar_arbiters_next_3_1_sva);
  assign mux_tmp_211 = MUX_s_1_2_2(or_tmp_253, mux_210_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign and_869_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_1_sva;
  assign nand_62_cse = ~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]) & Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1);
  assign or_974_nl = and_869_cse | Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 |
      or_tmp_253;
  assign mux_212_nl = MUX_s_1_2_2(mux_tmp_211, or_974_nl, Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1);
  assign or_972_nl = Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 | (~(nand_62_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 & (~ or_tmp_253)));
  assign mux_213_nl = MUX_s_1_2_2(mux_212_nl, or_972_nl, weight_mem_read_arbxbar_arbiters_next_3_3_sva);
  assign mux_214_nl = MUX_s_1_2_2(mux_tmp_211, mux_213_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign or_971_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3])
      | or_tmp_253;
  assign mux_208_nl = MUX_s_1_2_2(or_tmp_253, or_971_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign or_969_nl = weight_mem_read_arbxbar_arbiters_next_3_3_sva | and_869_cse
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]) | or_tmp_253;
  assign mux_209_nl = MUX_s_1_2_2(mux_208_nl, or_969_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign mux_tmp_215 = MUX_s_1_2_2(mux_214_nl, mux_209_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_873_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  assign and_875_cse = weight_mem_read_arbxbar_arbiters_next_3_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign or_tmp_265 = and_873_cse | and_869_cse | and_875_cse | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  assign mux_217_nl = MUX_s_1_2_2(or_tmp_265, mux_tmp_215, while_stage_0_5);
  assign nor_417_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_5_sva | (~ or_tmp_265));
  assign nor_418_nl = ~(while_mux_1445_tmp | (~ mux_tmp_215));
  assign mux_216_nl = MUX_s_1_2_2(nor_417_nl, nor_418_nl, while_stage_0_5);
  assign mux_218_nl = MUX_s_1_2_2(mux_217_nl, mux_216_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign and_dcpl_711 = mux_218_nl & (~(weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp));
  assign and_dcpl_713 = ~(weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign or_tmp_268 = and_873_cse | and_867_cse;
  assign or_tmp_270 = (Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]))
      | and_867_cse;
  assign or_986_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva | or_tmp_268;
  assign or_985_nl = Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 | or_tmp_270;
  assign mux_219_nl = MUX_s_1_2_2(or_986_nl, or_985_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign or_983_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3])
      | weight_mem_read_arbxbar_arbiters_next_3_1_sva | or_tmp_268;
  assign mux_tmp_220 = MUX_s_1_2_2(mux_219_nl, or_983_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_275 = and_873_cse | and_875_cse;
  assign mux_224_nl = MUX_s_1_2_2(or_tmp_268, or_tmp_270, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign or_994_nl = (Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_82_cse
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])) | and_867_cse;
  assign mux_tmp_225 = MUX_s_1_2_2(mux_224_nl, or_994_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign nor_423_cse = ~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]));
  assign mux_227_nl = MUX_s_1_2_2(or_tmp_275, mux_tmp_225, while_stage_0_5);
  assign nor_425_nl = ~(nor_423_cse | mux_227_nl);
  assign nor_426_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_5_sva | or_tmp_275);
  assign nor_427_nl = ~(while_mux_1445_tmp | mux_tmp_225);
  assign mux_226_nl = MUX_s_1_2_2(nor_426_nl, nor_427_nl, while_stage_0_5);
  assign mux_228_nl = MUX_s_1_2_2(nor_425_nl, mux_226_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign or_992_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva | or_tmp_275;
  assign mux_222_nl = MUX_s_1_2_2(or_992_nl, mux_tmp_220, while_stage_0_5);
  assign nor_428_nl = ~(nor_423_cse | mux_222_nl);
  assign nor_429_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_5_sva | weight_mem_read_arbxbar_arbiters_next_3_1_sva
      | or_tmp_275);
  assign nor_430_nl = ~(while_mux_1445_tmp | mux_tmp_220);
  assign mux_221_nl = MUX_s_1_2_2(nor_429_nl, nor_430_nl, while_stage_0_5);
  assign mux_223_nl = MUX_s_1_2_2(nor_428_nl, mux_221_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign mux_229_nl = MUX_s_1_2_2(mux_228_nl, mux_223_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign and_dcpl_714 = mux_229_nl & and_dcpl_713;
  assign or_1006_nl = nor_tmp_136 | and_867_cse;
  assign nand_16_nl = ~(nor_tmp_135 & (~ and_867_cse));
  assign mux_232_nl = MUX_s_1_2_2(or_1006_nl, nand_16_nl, weight_mem_read_arbxbar_arbiters_next_3_1_sva);
  assign mux_tmp_233 = MUX_s_1_2_2(and_867_cse, mux_232_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign or_1005_nl = and_869_cse | Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1
      | and_867_cse;
  assign mux_234_nl = MUX_s_1_2_2(mux_tmp_233, or_1005_nl, Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1);
  assign or_1003_nl = Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 | (~(nand_62_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 & (~ and_867_cse)));
  assign mux_235_nl = MUX_s_1_2_2(mux_234_nl, or_1003_nl, weight_mem_read_arbxbar_arbiters_next_3_3_sva);
  assign mux_236_nl = MUX_s_1_2_2(mux_tmp_233, mux_235_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign or_1002_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3])
      | and_867_cse;
  assign mux_230_nl = MUX_s_1_2_2(and_867_cse, or_1002_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign or_1000_nl = weight_mem_read_arbxbar_arbiters_next_3_3_sva | and_869_cse
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]) | and_867_cse;
  assign mux_231_nl = MUX_s_1_2_2(mux_230_nl, or_1000_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign mux_tmp_237 = MUX_s_1_2_2(mux_236_nl, mux_231_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_294 = and_873_cse | and_869_cse | and_875_cse;
  assign mux_tmp_238 = MUX_s_1_2_2(or_tmp_294, mux_tmp_237, while_stage_0_5);
  assign and_dcpl_721 = ~(mux_tmp_238 | weight_mem_read_arbxbar_xbar_1_for_3_4_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]));
  assign and_890_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  assign or_tmp_298 = and_890_cse | (weight_mem_read_arbxbar_arbiters_next_2_5_sva
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]));
  assign or_1011_nl = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign mux_tmp_241 = MUX_s_1_2_2(or_tmp_298, or_1011_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign nor_tmp_159 = Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign and_893_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) & Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1;
  assign or_tmp_300 = and_893_cse | nor_tmp_159;
  assign mux_tmp_242 = MUX_s_1_2_2(or_tmp_298, or_tmp_300, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign mux_245_nl = MUX_s_1_2_2(mux_tmp_242, mux_tmp_241, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_246_nl = MUX_s_1_2_2(or_tmp_298, mux_245_nl, while_stage_0_5);
  assign or_1016_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1
      | or_tmp_298;
  assign or_1015_nl = Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 | mux_tmp_242;
  assign or_1013_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1
      | mux_tmp_241;
  assign mux_243_nl = MUX_s_1_2_2(or_1015_nl, or_1013_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_244_nl = MUX_s_1_2_2(or_1016_nl, mux_243_nl, while_stage_0_5);
  assign mux_tmp_247 = MUX_s_1_2_2(mux_246_nl, mux_244_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign and_898_cse = weight_mem_read_arbxbar_arbiters_next_2_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign and_897_cse = weight_mem_read_arbxbar_arbiters_next_2_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign and_899_cse = weight_mem_read_arbxbar_arbiters_next_2_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign nand_17_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      & (~ or_tmp_298));
  assign mux_248_nl = MUX_s_1_2_2(nand_17_nl, or_tmp_298, and_897_cse);
  assign mux_249_nl = MUX_s_1_2_2(mux_248_nl, or_tmp_298, and_898_cse);
  assign mux_tmp_250 = MUX_s_1_2_2(mux_249_nl, or_tmp_298, and_899_cse);
  assign and_900_cse = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign or_tmp_307 = and_900_cse | mux_tmp_250;
  assign and_905_cse = Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign and_907_cse = Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign and_906_cse = Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign nand_18_nl = ~(Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      & (~ or_tmp_300));
  assign mux_252_nl = MUX_s_1_2_2(nand_18_nl, or_tmp_300, and_905_cse);
  assign mux_253_nl = MUX_s_1_2_2(mux_252_nl, or_tmp_300, and_906_cse);
  assign mux_254_nl = MUX_s_1_2_2(mux_253_nl, or_tmp_300, and_907_cse);
  assign mux_255_nl = MUX_s_1_2_2(mux_tmp_250, mux_254_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_1023_nl = (Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]))
      | mux_255_nl;
  assign or_1019_nl = and_900_cse | (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]))) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign mux_251_nl = MUX_s_1_2_2(or_tmp_307, or_1019_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign mux_256_nl = MUX_s_1_2_2(or_1023_nl, mux_251_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_257_itm = MUX_s_1_2_2(or_tmp_307, mux_256_nl, while_stage_0_5);
  assign or_1025_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign mux_258_nl = MUX_s_1_2_2((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]),
      or_1025_nl, weight_mem_read_arbxbar_arbiters_next_2_2_sva);
  assign mux_tmp_259 = MUX_s_1_2_2(and_898_cse, mux_258_nl, weight_mem_read_arbxbar_arbiters_next_2_5_sva);
  assign and_910_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  assign or_tmp_315 = and_910_cse | and_897_cse | and_899_cse | and_890_cse | mux_tmp_259;
  assign or_1024_nl = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign mux_tmp_260 = MUX_s_1_2_2(or_tmp_315, or_1024_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign or_tmp_317 = nor_tmp_159 | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign and_915_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) & Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1;
  assign or_1032_nl = and_893_cse | or_tmp_317;
  assign mux_261_nl = MUX_s_1_2_2(or_tmp_300, or_1032_nl, Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1);
  assign or_1035_nl = and_915_cse | and_905_cse | and_907_cse | mux_261_nl;
  assign mux_tmp_262 = MUX_s_1_2_2(or_tmp_315, or_1035_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_1037_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1
      | or_tmp_315;
  assign or_1036_nl = Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 | mux_tmp_262;
  assign or_1030_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1
      | mux_tmp_260;
  assign mux_263_nl = MUX_s_1_2_2(or_1036_nl, or_1030_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_264 = MUX_s_1_2_2(or_1037_nl, mux_263_nl, while_stage_0_5);
  assign mux_265_nl = MUX_s_1_2_2(mux_tmp_262, mux_tmp_260, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_266 = MUX_s_1_2_2(or_tmp_315, mux_265_nl, while_stage_0_5);
  assign or_1039_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])) |
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign mux_267_nl = MUX_s_1_2_2((~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])),
      or_1039_nl, weight_mem_read_arbxbar_arbiters_next_2_2_sva);
  assign or_1040_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva | mux_267_nl;
  assign or_1038_nl = weight_mem_read_arbxbar_arbiters_next_2_6_sva | mux_tmp_259;
  assign mux_268_nl = MUX_s_1_2_2(or_1040_nl, or_1038_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign or_tmp_329 = and_910_cse | and_897_cse | and_899_cse | mux_268_nl;
  assign or_1048_nl = Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]));
  assign or_1047_nl = Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 | nor_tmp_159;
  assign mux_270_nl = MUX_s_1_2_2(or_1048_nl, or_1047_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign or_1046_nl = Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]))
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign or_1045_nl = Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 | or_tmp_317;
  assign mux_269_nl = MUX_s_1_2_2(or_1046_nl, or_1045_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign mux_271_nl = MUX_s_1_2_2(mux_270_nl, mux_269_nl, Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1);
  assign or_1051_nl = and_915_cse | and_905_cse | and_907_cse | mux_271_nl;
  assign mux_272_nl = MUX_s_1_2_2(or_tmp_329, or_1051_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_1044_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2])
      | or_tmp_329;
  assign mux_273_nl = MUX_s_1_2_2(mux_272_nl, or_1044_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_274_nl = MUX_s_1_2_2(or_tmp_329, mux_273_nl, while_stage_0_5);
  assign mux_275_nl = MUX_s_1_2_2(mux_274_nl, mux_tmp_266, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]);
  assign mux_276_itm = MUX_s_1_2_2(mux_275_nl, mux_tmp_264, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign or_tmp_338 = and_899_cse | and_898_cse;
  assign or_1057_nl = weight_mem_read_arbxbar_arbiters_next_2_2_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]));
  assign or_1056_nl = weight_mem_read_arbxbar_arbiters_next_2_1_sva | and_898_cse;
  assign mux_277_nl = MUX_s_1_2_2(or_1057_nl, or_1056_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign or_1055_nl = weight_mem_read_arbxbar_arbiters_next_2_3_sva | or_tmp_338;
  assign mux_278_nl = MUX_s_1_2_2(mux_277_nl, or_1055_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign or_1054_nl = weight_mem_read_arbxbar_arbiters_next_2_4_sva | and_897_cse
      | or_tmp_338;
  assign mux_tmp_279 = MUX_s_1_2_2(mux_278_nl, or_1054_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign or_tmp_345 = and_907_cse | and_906_cse;
  assign or_1064_nl = Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]));
  assign or_1063_nl = Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 | and_906_cse;
  assign mux_280_nl = MUX_s_1_2_2(or_1064_nl, or_1063_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign or_1062_nl = Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 | or_tmp_345;
  assign mux_281_nl = MUX_s_1_2_2(mux_280_nl, or_1062_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign or_1061_nl = Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 | and_905_cse |
      or_tmp_345;
  assign mux_282_nl = MUX_s_1_2_2(mux_281_nl, or_1061_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign mux_283_nl = MUX_s_1_2_2(mux_tmp_279, mux_282_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign or_1058_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2])
      | mux_tmp_279;
  assign mux_284_nl = MUX_s_1_2_2(mux_283_nl, or_1058_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_285_nl = MUX_s_1_2_2(mux_tmp_279, mux_284_nl, while_stage_0_5);
  assign and_dcpl_725 = (~ mux_285_nl) & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]))) & and_dcpl_635;
  assign while_mux_1483_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_287_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      while_mux_1483_nl, while_stage_0_5);
  assign and_dcpl_726 = mux_287_nl & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign or_dcpl_715 = and_dcpl_726 | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign and_dcpl_727 = ~(weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp);
  assign nor_tmp_197 = while_mux_1429_cse_1 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign nor_tmp_199 = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign nand_20_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      & (~ nor_tmp_199));
  assign nand_19_nl = ~(while_mux_1435_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      & (~ nor_tmp_197));
  assign mux_288_nl = MUX_s_1_2_2(nand_20_nl, nand_19_nl, while_stage_0_5);
  assign or_1067_nl = weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  assign mux_289_nl = MUX_s_1_2_2(mux_288_nl, and_dcpl_726, or_1067_nl);
  assign and_dcpl_728 = (~ mux_289_nl) & and_dcpl_727;
  assign and_dcpl_731 = and_dcpl_727 & (~ weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp)
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp));
  assign not_tmp_456 = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]));
  assign or_tmp_353 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) | not_tmp_456;
  assign not_tmp_457 = ~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]));
  assign mux_291_nl = MUX_s_1_2_2(not_tmp_457, or_tmp_353, Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1);
  assign nor_442_nl = ~(and_1000_cse | mux_291_nl);
  assign mux_290_nl = MUX_s_1_2_2(not_tmp_457, or_tmp_353, while_mux_1429_cse_1);
  assign nor_443_nl = ~(and_1001_cse | mux_290_nl);
  assign mux_292_nl = MUX_s_1_2_2(nor_442_nl, nor_443_nl, while_stage_0_5);
  assign and_dcpl_732 = mux_292_nl & and_dcpl_731;
  assign mux_293_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_1_sva,
      while_mux_1435_tmp, while_stage_0_5);
  assign and_dcpl_738 = (~(mux_293_nl & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])))
      & not_tmp_456 & (~ (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])) &
      (~(weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp));
  assign and_937_cse = weight_mem_read_arbxbar_arbiters_next_0_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign and_936_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) & weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  assign or_tmp_360 = and_936_cse | and_937_cse;
  assign or_1076_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign mux_tmp_295 = MUX_s_1_2_2(or_tmp_360, or_1076_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign or_1079_cse = and_1007_cse | and_1008_cse;
  assign mux_tmp_296 = MUX_s_1_2_2(or_tmp_360, or_1079_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign mux_299_nl = MUX_s_1_2_2(mux_tmp_296, mux_tmp_295, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_300_nl = MUX_s_1_2_2(or_tmp_360, mux_299_nl, while_stage_0_5);
  assign or_1081_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | or_tmp_360;
  assign or_1080_nl = Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 | mux_tmp_296;
  assign or_1078_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | mux_tmp_295;
  assign mux_297_nl = MUX_s_1_2_2(or_1080_nl, or_1078_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_298_nl = MUX_s_1_2_2(or_1081_nl, mux_297_nl, while_stage_0_5);
  assign mux_tmp_301 = MUX_s_1_2_2(mux_300_nl, mux_298_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign and_944_cse = weight_mem_read_arbxbar_arbiters_next_0_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]);
  assign and_943_cse = weight_mem_read_arbxbar_arbiters_next_0_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign and_945_cse = weight_mem_read_arbxbar_arbiters_next_0_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign nand_21_nl = ~(weight_mem_read_arbxbar_arbiters_next_0_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      & (~ or_tmp_360));
  assign mux_302_nl = MUX_s_1_2_2(nand_21_nl, or_tmp_360, and_943_cse);
  assign mux_303_nl = MUX_s_1_2_2(mux_302_nl, or_tmp_360, and_944_cse);
  assign mux_tmp_304 = MUX_s_1_2_2(mux_303_nl, or_tmp_360, and_945_cse);
  assign or_tmp_369 = and_1009_cse | mux_tmp_304;
  assign nand_22_nl = ~(Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      & (~ or_1079_cse));
  assign mux_306_nl = MUX_s_1_2_2(nand_22_nl, or_1079_cse, and_1004_cse);
  assign mux_307_nl = MUX_s_1_2_2(mux_306_nl, or_1079_cse, and_1003_cse);
  assign mux_308_nl = MUX_s_1_2_2(mux_307_nl, or_1079_cse, and_1006_cse);
  assign mux_309_nl = MUX_s_1_2_2(mux_tmp_304, mux_308_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign or_1088_nl = and_1002_cse | mux_309_nl;
  assign or_1084_nl = and_1009_cse | (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]))) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign mux_305_nl = MUX_s_1_2_2(or_tmp_369, or_1084_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign mux_310_nl = MUX_s_1_2_2(or_1088_nl, mux_305_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_311_itm = MUX_s_1_2_2(or_tmp_369, mux_310_nl, while_stage_0_5);
  assign and_958_cse = weight_mem_read_arbxbar_arbiters_next_0_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign or_tmp_377 = and_944_cse | and_943_cse | and_958_cse | and_945_cse | and_936_cse
      | and_937_cse;
  assign or_1089_nl = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign mux_tmp_312 = MUX_s_1_2_2(or_tmp_377, or_1089_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign or_1104_nl = weight_mem_read_arbxbar_arbiters_next_0_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]));
  assign or_1103_nl = weight_mem_read_arbxbar_arbiters_next_0_5_sva | and_937_cse;
  assign mux_316_nl = MUX_s_1_2_2(or_1104_nl, or_1103_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign or_tmp_391 = and_944_cse | and_943_cse | and_958_cse | and_945_cse | mux_316_nl;
  assign mux_tmp_320 = MUX_s_1_2_2(or_tmp_391, or_tmp_377, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign or_1111_nl = Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]));
  assign or_1110_nl = Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 | and_1008_cse;
  assign mux_318_nl = MUX_s_1_2_2(or_1111_nl, or_1110_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign or_1115_nl = and_1003_cse | and_1004_cse | and_1005_cse | and_1006_cse |
      mux_318_nl;
  assign mux_319_nl = MUX_s_1_2_2(or_1115_nl, or_1140_cse, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign mux_321_nl = MUX_s_1_2_2(mux_tmp_320, mux_319_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign or_1109_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0])
      | or_tmp_391;
  assign mux_317_nl = MUX_s_1_2_2(or_1109_nl, mux_tmp_312, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign mux_322_nl = MUX_s_1_2_2(mux_321_nl, mux_317_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_323_nl = MUX_s_1_2_2(mux_tmp_320, mux_322_nl, while_stage_0_5);
  assign or_1102_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | or_tmp_377;
  assign or_1101_nl = Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 | mux_335_cse;
  assign or_1095_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | mux_tmp_312;
  assign mux_314_nl = MUX_s_1_2_2(or_1101_nl, or_1095_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_315_nl = MUX_s_1_2_2(or_1102_nl, mux_314_nl, while_stage_0_5);
  assign mux_324_itm = MUX_s_1_2_2(mux_323_nl, mux_315_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign or_tmp_399 = and_943_cse | and_944_cse;
  assign or_1121_nl = weight_mem_read_arbxbar_arbiters_next_0_1_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]));
  assign or_1120_nl = weight_mem_read_arbxbar_arbiters_next_0_2_sva | and_944_cse;
  assign mux_325_nl = MUX_s_1_2_2(or_1121_nl, or_1120_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign or_1119_nl = weight_mem_read_arbxbar_arbiters_next_0_3_sva | or_tmp_399;
  assign mux_326_nl = MUX_s_1_2_2(mux_325_nl, or_1119_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign or_1118_nl = weight_mem_read_arbxbar_arbiters_next_0_4_sva | and_958_cse
      | or_tmp_399;
  assign mux_tmp_327 = MUX_s_1_2_2(mux_326_nl, or_1118_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign or_tmp_406 = and_1004_cse | and_1003_cse;
  assign or_1128_nl = Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]));
  assign or_1127_nl = Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 | and_1003_cse;
  assign mux_328_nl = MUX_s_1_2_2(or_1128_nl, or_1127_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign or_1126_nl = Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 | or_tmp_406;
  assign mux_329_nl = MUX_s_1_2_2(mux_328_nl, or_1126_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign or_1125_nl = Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 | and_1005_cse |
      or_tmp_406;
  assign mux_330_nl = MUX_s_1_2_2(mux_329_nl, or_1125_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign mux_331_nl = MUX_s_1_2_2(mux_tmp_327, mux_330_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign or_1122_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0])
      | mux_tmp_327;
  assign mux_332_nl = MUX_s_1_2_2(mux_331_nl, or_1122_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_333_nl = MUX_s_1_2_2(mux_tmp_327, mux_332_nl, while_stage_0_5);
  assign and_dcpl_742 = (~ mux_333_nl) & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]))) & and_dcpl_621;
  assign or_tmp_418 = and_1009_cse | or_tmp_377;
  assign or_dcpl_717 = ~(weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign and_580_nl = fsm_output & (~ weight_mem_run_3_for_land_4_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
      weight_port_read_out_data_3_15_sva_dfm_1, and_580_nl);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[255:240];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_c = weight_mem_run_3_for_5_mux_62_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[239:224];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_a = weight_port_read_out_data_7_1_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_b = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[31:16];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_c = weight_port_read_out_data_7_0_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_1_d = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[15:0];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_2_a = weight_port_read_out_data_7_3_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_2_b = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[63:48];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_2_c = weight_port_read_out_data_7_2_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_2_d = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[47:32];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_3_a = weight_port_read_out_data_7_5_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_3_b = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[95:80];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_3_c = weight_port_read_out_data_7_4_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_3_d = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[79:64];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_4_a = weight_port_read_out_data_7_7_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_4_b = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[127:112];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_4_c = weight_port_read_out_data_7_6_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_4_d = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[111:96];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_5_a = weight_port_read_out_data_7_9_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_5_b = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[159:144];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_5_c = weight_port_read_out_data_7_8_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_5_d = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[143:128];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_6_a = weight_port_read_out_data_7_11_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_6_b = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[191:176];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_6_c = weight_port_read_out_data_7_10_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_6_d = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[175:160];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_7_a = weight_port_read_out_data_7_13_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_7_b = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[223:208];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_7_c = weight_port_read_out_data_7_12_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_7_d = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[207:192];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_8_a = weight_port_read_out_data_7_15_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[255:240];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_8_c = weight_port_read_out_data_7_14_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[239:224];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_9_a = {weight_port_read_out_data_0_1_sva_dfm_1_1_15
      , weight_port_read_out_data_0_1_sva_dfm_1_1_14_0};
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[31:16];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_9_c = weight_port_read_out_data_0_0_sva_dfm_1_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[15:0];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_10_a = weight_port_read_out_data_0_3_sva_dfm_1_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[63:48];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_10_c = weight_port_read_out_data_0_2_sva_dfm_1_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[47:32];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_11_a = weight_mem_run_3_for_5_mux_5_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[95:80];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_11_c = weight_mem_run_3_for_5_mux_4_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[79:64];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_12_a = weight_mem_run_3_for_5_mux_7_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[127:112];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_12_c = weight_mem_run_3_for_5_mux_6_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[111:96];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_13_a = weight_mem_run_3_for_5_mux_9_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[159:144];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_13_c = weight_mem_run_3_for_5_mux_8_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[143:128];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_14_a = rva_out_reg_data_95_80_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[191:176];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_14_c = rva_out_reg_data_111_96_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[175:160];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_15_a = weight_mem_run_3_for_5_mux_13_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[223:208];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_15_c = weight_mem_run_3_for_5_mux_12_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5[207:192];
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_16_a = weight_mem_run_3_for_5_mux_15_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_16_c = weight_mem_run_3_for_5_mux_14_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_17_a = weight_mem_run_3_for_5_mux_97_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_17_c = weight_mem_run_3_for_5_mux_96_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_18_a = weight_mem_run_3_for_5_mux_99_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_18_c = weight_mem_run_3_for_5_mux_98_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_19_a = rva_out_reg_data_143_128_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_19_c = rva_out_reg_data_127_112_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_20_a = rva_out_reg_data_175_160_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_20_c = rva_out_reg_data_159_144_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_21_a = rva_out_reg_data_207_192_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_21_c = rva_out_reg_data_191_176_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_22_a = rva_out_reg_data_239_224_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_22_c = rva_out_reg_data_223_208_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_23_a = rva_out_reg_data_79_64_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_23_c = rva_out_reg_data_255_240_sva_dfm_4_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_24_a = weight_mem_run_3_for_5_mux_111_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_24_c = weight_mem_run_3_for_5_mux_110_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_25_a = weight_mem_run_3_for_5_mux_17_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_25_c = weight_mem_run_3_for_5_mux_16_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_26_a = weight_mem_run_3_for_5_mux_19_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_26_c = weight_mem_run_3_for_5_mux_18_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_27_a = weight_mem_run_3_for_5_mux_21_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_27_c = weight_mem_run_3_for_5_mux_20_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_28_a = weight_mem_run_3_for_5_mux_23_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_28_c = weight_mem_run_3_for_5_mux_22_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_29_a = weight_mem_run_3_for_5_mux_25_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_29_c = weight_mem_run_3_for_5_mux_24_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_30_a = weight_mem_run_3_for_5_mux_27_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_30_c = weight_mem_run_3_for_5_mux_26_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_31_a = weight_mem_run_3_for_5_mux_29_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_31_c = weight_mem_run_3_for_5_mux_28_itm_1;
  assign and_579_nl = fsm_output & (~ weight_mem_run_3_for_land_2_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_32_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
      weight_port_read_out_data_1_15_sva_dfm_1, and_579_nl);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_32_c = weight_mem_run_3_for_5_mux_30_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_33_a = weight_mem_run_3_for_5_mux_81_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_33_c = weight_mem_run_3_for_5_mux_80_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_34_a = weight_mem_run_3_for_5_mux_83_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_34_c = weight_mem_run_3_for_5_mux_82_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_35_a = weight_mem_run_3_for_5_mux_85_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_35_c = weight_mem_run_3_for_5_mux_84_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_36_a = weight_mem_run_3_for_5_mux_87_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_36_c = weight_mem_run_3_for_5_mux_86_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_37_a = weight_mem_run_3_for_5_mux_89_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_37_c = weight_mem_run_3_for_5_mux_88_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_38_a = weight_mem_run_3_for_5_mux_91_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_38_c = weight_mem_run_3_for_5_mux_90_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_39_a = weight_mem_run_3_for_5_mux_93_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_39_c = weight_mem_run_3_for_5_mux_92_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_40_a = weight_port_read_out_data_5_15_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_40_c = weight_port_read_out_data_5_14_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_41_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
      weight_port_read_out_data_2_1_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_41_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001,
      weight_port_read_out_data_2_0_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_42_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002,
      weight_port_read_out_data_2_3_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_42_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003,
      weight_port_read_out_data_2_2_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_43_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004,
      weight_port_read_out_data_2_5_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_43_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005,
      weight_port_read_out_data_2_4_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_44_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006,
      weight_port_read_out_data_2_7_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_44_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007,
      weight_port_read_out_data_2_6_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_45_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008,
      weight_port_read_out_data_2_9_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_45_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009,
      weight_port_read_out_data_2_8_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_46_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010,
      weight_port_read_out_data_2_11_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_46_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011,
      weight_port_read_out_data_2_10_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_47_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012,
      weight_port_read_out_data_2_13_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_47_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013,
      weight_port_read_out_data_2_12_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_48_a = weight_mem_run_3_for_5_mux_47_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_48_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014,
      weight_port_read_out_data_2_14_sva_dfm_1, and_dcpl_568);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_49_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
      weight_port_read_out_data_4_1_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_49_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001,
      weight_port_read_out_data_4_0_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_50_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002,
      weight_port_read_out_data_4_3_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_50_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003,
      weight_port_read_out_data_4_2_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_51_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004,
      weight_port_read_out_data_4_5_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_51_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005,
      weight_port_read_out_data_4_4_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_52_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006,
      weight_port_read_out_data_4_7_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_52_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007,
      weight_port_read_out_data_4_6_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_53_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008,
      weight_port_read_out_data_4_9_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_53_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009,
      weight_port_read_out_data_4_8_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_54_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010,
      weight_port_read_out_data_4_11_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_54_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011,
      weight_port_read_out_data_4_10_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_55_a = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012,
      weight_port_read_out_data_4_13_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_55_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013,
      weight_port_read_out_data_4_12_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_56_a = weight_mem_run_3_for_5_mux_79_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_56_c = MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014,
      weight_port_read_out_data_4_14_sva_dfm_1, and_dcpl_567);
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_57_a = weight_mem_run_3_for_5_mux_49_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_57_c = weight_mem_run_3_for_5_mux_48_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_58_a = weight_mem_run_3_for_5_mux_51_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_58_c = weight_mem_run_3_for_5_mux_50_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_59_a = weight_mem_run_3_for_5_mux_53_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_59_c = weight_mem_run_3_for_5_mux_52_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_60_a = weight_mem_run_3_for_5_mux_55_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_60_c = weight_mem_run_3_for_5_mux_54_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_61_a = weight_mem_run_3_for_5_mux_57_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_61_c = weight_mem_run_3_for_5_mux_56_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_62_a = weight_mem_run_3_for_5_mux_59_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_62_c = weight_mem_run_3_for_5_mux_58_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_63_a = weight_mem_run_3_for_5_mux_61_itm_1;
  assign Datapath_for_4_ProductSum_for_acc_9_cmp_63_c = weight_mem_run_3_for_5_mux_60_itm_1;
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0));
  assign weight_mem_banks_write_if_for_if_and_35_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_36_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_37_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_38_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_39_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_40_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_41_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      , weight_mem_banks_write_if_for_if_and_35_nl , weight_mem_banks_write_if_for_if_and_36_nl
      , weight_mem_banks_write_if_for_if_and_37_nl , weight_mem_banks_write_if_for_if_and_38_nl
      , weight_mem_banks_write_if_for_if_and_39_nl , weight_mem_banks_write_if_for_if_and_40_nl
      , weight_mem_banks_write_if_for_if_and_41_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0});
  assign weight_mem_banks_write_if_for_if_mux_7_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      , weight_mem_banks_write_if_for_if_mux_7_nl};
  assign nor_461_nl = ~((~ PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3) |
      PECore_RunFSM_switch_lp_equal_tmp_1_2);
  assign mux_123_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_461_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff = mux_123_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_2[14:3];
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff = and_dcpl_154;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0));
  assign weight_mem_banks_write_if_for_if_and_28_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_29_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_30_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_31_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_32_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_33_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_34_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      , weight_mem_banks_write_if_for_if_and_28_nl , weight_mem_banks_write_if_for_if_and_29_nl
      , weight_mem_banks_write_if_for_if_and_30_nl , weight_mem_banks_write_if_for_if_and_31_nl
      , weight_mem_banks_write_if_for_if_and_32_nl , weight_mem_banks_write_if_for_if_and_33_nl
      , weight_mem_banks_write_if_for_if_and_34_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0});
  assign weight_mem_banks_write_if_for_if_mux_6_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      , weight_mem_banks_write_if_for_if_mux_6_nl};
  assign nor_460_nl = ~(PECore_UpdateFSM_switch_lp_equal_tmp_2_3 | (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_122_nl = MUX_s_1_2_2(or_tmp_111, nor_460_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff = mux_122_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff = and_dcpl_156;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0));
  assign weight_mem_banks_write_if_for_if_and_21_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_22_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_23_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_24_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_25_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_26_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_27_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      , weight_mem_banks_write_if_for_if_and_21_nl , weight_mem_banks_write_if_for_if_and_22_nl
      , weight_mem_banks_write_if_for_if_and_23_nl , weight_mem_banks_write_if_for_if_and_24_nl
      , weight_mem_banks_write_if_for_if_and_25_nl , weight_mem_banks_write_if_for_if_and_26_nl
      , weight_mem_banks_write_if_for_if_and_27_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0});
  assign weight_mem_banks_write_if_for_if_mux_5_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      , weight_mem_banks_write_if_for_if_mux_5_nl};
  assign nor_459_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_3) | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]));
  assign mux_121_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_459_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff = mux_121_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff = and_dcpl_158;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0));
  assign weight_mem_banks_write_if_for_if_and_14_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_15_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_16_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_17_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_18_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_19_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_20_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      , weight_mem_banks_write_if_for_if_and_14_nl , weight_mem_banks_write_if_for_if_and_15_nl
      , weight_mem_banks_write_if_for_if_and_16_nl , weight_mem_banks_write_if_for_if_and_17_nl
      , weight_mem_banks_write_if_for_if_and_18_nl , weight_mem_banks_write_if_for_if_and_19_nl
      , weight_mem_banks_write_if_for_if_and_20_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0});
  assign weight_mem_banks_write_if_for_if_mux_4_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      , weight_mem_banks_write_if_for_if_mux_4_nl};
  assign nor_458_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3) | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]));
  assign mux_120_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_458_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff = mux_120_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff = and_dcpl_160;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0));
  assign weight_mem_banks_write_if_for_if_and_7_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_9_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_10_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_11_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_12_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_13_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      , weight_mem_banks_write_if_for_if_and_7_nl , weight_mem_banks_write_if_for_if_and_8_nl
      , weight_mem_banks_write_if_for_if_and_9_nl , weight_mem_banks_write_if_for_if_and_10_nl
      , weight_mem_banks_write_if_for_if_and_11_nl , weight_mem_banks_write_if_for_if_and_12_nl
      , weight_mem_banks_write_if_for_if_and_13_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0});
  assign weight_mem_banks_write_if_for_if_mux_3_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      , weight_mem_banks_write_if_for_if_mux_3_nl};
  assign nor_457_nl = ~((~ pe_manager_base_weight_slc_pe_manager_base_weight_2_0_380_itm_1)
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]));
  assign mux_119_nl = MUX_s_1_2_2(or_50_cse, nor_457_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff = mux_119_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff = and_dcpl_162;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_14_lpi_1_dfm_1_2_6 , weight_write_data_data_0_13_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_12_lpi_1_dfm_1_2_6 , weight_write_data_data_0_11_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_10_lpi_1_dfm_1_2_6 , weight_write_data_data_0_9_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_8_lpi_1_dfm_1_2_6 , weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0));
  assign weight_mem_banks_write_if_for_if_and_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_1_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_2_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_3_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_5_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl ,
      weight_mem_banks_write_if_for_if_and_nl , weight_mem_banks_write_if_for_if_and_1_nl
      , weight_mem_banks_write_if_for_if_and_2_nl , weight_mem_banks_write_if_for_if_and_3_nl
      , weight_mem_banks_write_if_for_if_and_4_nl , weight_mem_banks_write_if_for_if_and_5_nl
      , weight_mem_banks_write_if_for_if_and_6_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0});
  assign weight_mem_banks_write_if_for_if_mux_2_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      , weight_mem_banks_write_if_for_if_mux_2_nl};
  assign nor_456_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1)
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]));
  assign mux_118_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_456_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff = mux_118_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff = and_dcpl_164;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_14_lpi_1_dfm_1_3_2 , weight_write_data_data_0_13_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_12_lpi_1_dfm_1_3_2 , weight_write_data_data_0_11_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_10_lpi_1_dfm_1_3_2 , weight_write_data_data_0_9_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_8_lpi_1_dfm_1_3_2 , weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_1_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_54_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0,
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_1_nl
      , weight_mem_banks_write_if_for_if_mux_54_nl};
  assign nor_455_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_1);
  assign mux_117_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_455_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff = mux_117_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_3_14_3;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff = and_dcpl_546;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d = {weight_write_data_data_0_15_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_14_lpi_1_dfm_1_3_2 , weight_write_data_data_0_13_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_12_lpi_1_dfm_1_3_2 , weight_write_data_data_0_11_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_10_lpi_1_dfm_1_3_2 , weight_write_data_data_0_9_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_8_lpi_1_dfm_1_3_2 , weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_53_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0,
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_nl
      , weight_mem_banks_write_if_for_if_mux_53_nl};
  assign nor_454_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1);
  assign mux_116_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_454_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff = mux_116_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff = and_dcpl_544;
  assign and_dcpl_743 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1
      & (weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[1]);
  assign or_dcpl = and_dcpl_743 | ((weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_itm_1);
  assign or_dcpl_719 = (nor_335_cse & (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]))
      | ((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]) & (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]))
      | (and_dcpl_657 & (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]));
  assign or_dcpl_720 = and_dcpl_743 | ((weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_231_itm_1);
  assign or_197_nl = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      | not_tmp_139;
  assign mux_44_nl = MUX_s_1_2_2((~ or_tmp_35), or_197_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1);
  assign weight_mem_banks_load_store_for_else_and_80_ssc = PECoreRun_wen & mux_44_nl
      & and_dcpl_56;
  assign weight_port_read_out_data_and_209_enex5 = weight_port_read_out_data_and_170_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_298_enex5 = rva_out_reg_data_and_128_cse & reg_rva_out_reg_data_30_25_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_299_enex5 = rva_out_reg_data_and_166_cse & reg_rva_out_reg_data_30_25_sva_dfm_2_enexo;
  assign nor_340_nl = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2) | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1
      | input_read_req_valid_lpi_1_dfm_1_3 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 | PECore_DecodeAxiRead_switch_lp_nor_tmp_3
      | rva_in_reg_rw_sva_3 | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_363_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1);
  assign mux_68_nl = MUX_s_1_2_2(mux_tmp_51, nor_340_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign rva_out_reg_data_and_168_ssc = PECoreRun_wen & mux_68_nl & while_stage_0_5;
  assign rva_out_reg_data_and_300_enex5 = rva_out_reg_data_and_168_ssc & reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  assign accum_vector_data_and_16_cse = and_dcpl_24 & fsm_output;
  assign weight_mem_run_3_for_5_and_158_ssc = reg_weight_mem_run_3_for_5_and_146_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_159_ssc = reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_160_ssc = reg_weight_mem_run_3_for_5_and_148_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_161_ssc = reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_164_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_port_read_out_data_and_128_ssc = PECoreRun_wen & and_dcpl_45;
  assign weight_port_read_out_data_and_210_enex5 = weight_port_read_out_data_and_164_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_301_enex5 = rva_out_reg_data_and_68_cse & reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  assign weight_port_read_out_data_and_211_enex5 = weight_port_read_out_data_and_166_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo;
  assign rva_out_reg_data_and_89_ssc = PECoreRun_wen & and_dcpl_348 & (~ rva_in_reg_rw_sva_st_1_7)
      & (~(rva_in_reg_rw_sva_st_7 | PECore_DecodeAxiRead_switch_lp_nor_tmp_7 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7))
      & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & while_stage_0_9 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5
      | input_read_req_valid_lpi_1_dfm_1_7));
  assign rva_out_reg_data_and_302_enex5 = rva_out_reg_data_and_89_ssc & reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_130_ssc = PECoreRun_wen & and_dcpl_195 & (~(rva_in_reg_rw_sva_5
      & rva_in_reg_rw_sva_st_1_5));
  assign weight_port_read_out_data_0_1_sva_mx0_15 = MUX1HOT_s_1_3_2(weight_port_read_out_data_0_1_sva_dfm_1_15,
      weight_port_read_out_data_0_1_sva_dfm_1_1_15, weight_port_read_out_data_0_1_sva_15,
      {and_dcpl_367 , and_dcpl_320 , (~ while_stage_0_8)});
  assign weight_port_read_out_data_0_1_sva_mx0_14_0 = MUX1HOT_v_15_3_2(weight_port_read_out_data_0_1_sva_dfm_1_14_0,
      weight_port_read_out_data_0_1_sva_dfm_1_1_14_0, weight_port_read_out_data_0_1_sva_14_0,
      {and_dcpl_367 , and_dcpl_320 , (~ while_stage_0_8)});
  assign rva_out_reg_data_35_32_sva_dfm_6_mx1_3_2 = MUX_v_2_2_2(rva_out_reg_data_35_32_sva_dfm_4_1_3_2,
      rva_out_reg_data_35_32_sva_dfm_6_rsp_0, or_dcpl_706);
  assign rva_out_reg_data_35_32_sva_dfm_6_mx1_1_0 = MUX_v_2_2_2(rva_out_reg_data_35_32_sva_dfm_4_1_1_0,
      rva_out_reg_data_35_32_sva_dfm_6_rsp_1, or_dcpl_706);
  assign rva_out_reg_data_and_303_enex5 = rva_out_reg_data_and_26_cse & reg_rva_out_reg_data_30_25_sva_dfm_8_enexo;
  assign and_dcpl_808 = fsm_output & while_stage_0_7;
  assign or_dcpl_752 = weight_mem_run_3_for_5_and_142_itm_1 | weight_mem_run_3_for_5_and_140_itm_2;
  assign or_dcpl_753 = weight_mem_run_3_for_5_and_144_itm_1 | weight_mem_run_3_for_5_and_143_itm_1;
  assign or_dcpl_761 = weight_mem_run_3_for_5_and_135_itm_2 | weight_mem_run_3_for_5_and_126_itm_2;
  assign or_dcpl_766 = weight_mem_run_3_for_5_and_144_itm_1 | weight_mem_run_3_for_5_and_135_itm_2;
  assign or_dcpl_774 = weight_mem_run_3_for_5_and_126_itm_2 | weight_mem_run_3_for_5_and_140_itm_2;
  assign or_dcpl_792 = weight_mem_run_3_for_5_and_143_itm_1 | weight_mem_run_3_for_5_and_126_itm_2;
  assign or_tmp_441 = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  assign or_1312_nl = rva_in_PopNB_mioi_return_rsc_z_mxwt | (state_2_1_sva[1]) |
      (~((state_2_1_sva[0]) & state_0_sva & reg_rva_in_PopNB_mioi_iswt0_cse));
  assign or_1310_nl = PECore_UpdateFSM_switch_lp_equal_tmp_3_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1);
  assign mux_381_nl = MUX_s_1_2_2(or_1312_nl, or_1310_nl, while_stage_0_3);
  assign or_1308_nl = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  assign mux_382_nl = MUX_s_1_2_2(mux_381_nl, or_1308_nl, while_stage_0_4);
  assign or_1307_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_3 | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_3);
  assign mux_383_nl = MUX_s_1_2_2(mux_382_nl, or_1307_nl, while_stage_0_5);
  assign or_1305_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse);
  assign mux_384_nl = MUX_s_1_2_2(mux_383_nl, or_1305_nl, while_stage_0_6);
  assign or_1303_nl = PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_5);
  assign mux_385_nl = MUX_s_1_2_2(mux_384_nl, or_1303_nl, while_stage_0_7);
  assign or_1301_nl = PECore_RunMac_PECore_RunMac_if_and_svs_st_6 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_6);
  assign mux_386_nl = MUX_s_1_2_2(mux_385_nl, or_1301_nl, while_stage_0_8);
  assign or_1299_nl = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_7) | PECore_RunMac_PECore_RunMac_if_and_svs_st_7
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  assign mux_387_nl = MUX_s_1_2_2(mux_386_nl, or_1299_nl, while_stage_0_9);
  assign or_1298_nl = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_8) | PECore_RunMac_PECore_RunMac_if_and_svs_st_8
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  assign mux_388_nl = MUX_s_1_2_2(mux_387_nl, or_1298_nl, while_stage_0_10);
  assign or_1297_nl = (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_9) | PECore_RunMac_PECore_RunMac_if_and_svs_st_9
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9;
  assign mux_tmp_376 = MUX_s_1_2_2(mux_388_nl, or_1297_nl, while_stage_0_11);
  assign and_1120_tmp = (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | (~ while_stage_0_11)
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_8 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9)
      & while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen;
  assign data_in_tmp_operator_2_for_and_tmp = PECoreRun_wen & and_dcpl_45 & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign data_in_tmp_operator_2_for_and_31_tmp = PECoreRun_wen & and_dcpl_45 & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign rva_in_reg_data_and_tmp = PECoreRun_wen & and_dcpl_282 & (and_279_cse |
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign input_mem_banks_read_1_read_data_and_4_tmp = PECoreRun_wen & (and_352_cse
      | ((~ reg_rva_in_reg_rw_sva_st_1_1_cse) & input_read_req_valid_lpi_1_dfm_1_1
      & and_dcpl_172));
  assign nand_36_nl = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign nor_nl = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5));
  assign mux_nl = MUX_s_1_2_2(nand_36_nl, nor_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_5);
  assign mux_1_nl = MUX_s_1_2_2(mux_nl, or_tmp, rva_in_reg_rw_sva_st_1_5);
  assign weight_port_read_out_data_and_127_tmp = PECoreRun_wen & (~ mux_1_nl) & while_stage_0_7;
  assign input_mem_banks_read_read_data_and_54_tmp = PECoreRun_wen & (~((~((~ rva_in_reg_rw_sva_st_1_4)
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)))
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
      & while_stage_0_6;
  assign pe_manager_base_input_and_tmp = PECoreRun_wen & ((nand_83_cse & while_stage_0_3)
      | and_dcpl_180);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_63_cse <= 1'b0;
      reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_40_cse <= 1'b0;
      reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_7_cse <= 1'b0;
      reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_1_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_act_port_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      pe_config_manager_counter_sva_dfm_3_1 <= 4'b0000;
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= 1'b0;
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= 1'b0;
      while_stage_0_3 <= 1'b0;
      while_stage_0_4 <= 1'b0;
      while_stage_0_5 <= 1'b0;
      while_stage_0_6 <= 1'b0;
      while_stage_0_7 <= 1'b0;
      while_stage_0_8 <= 1'b0;
      while_stage_0_9 <= 1'b0;
      while_stage_0_10 <= 1'b0;
      while_stage_0_11 <= 1'b0;
      while_stage_0_12 <= 1'b0;
      while_stage_0_13 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_359_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_153_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_141_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_5_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_4_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_1 <= 1'b0;
      input_read_addrs_sva_1_1 <= 8'b00000000;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= 1'b0;
      weight_port_read_out_data_0_1_sva_15 <= 1'b0;
    end
    else if ( PECoreRun_wen ) begin
      reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_63_cse <= and_535_rmff;
      reg_Datapath_for_4_ProductSum_for_acc_9_cmp_cgo_ir_40_cse <= and_538_rmff;
      reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_7_cse <= and_541_rmff;
      reg_PECore_RunScale_if_for_1_scaled_val_mul_1_cmp_cgo_ir_1_cse <= and_544_rmff;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= and_548_rmff;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= and_551_rmff;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= and_555_rmff;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= and_558_rmff;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= and_561_rmff;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= and_564_rmff;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= and_567_rmff;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= and_570_rmff;
      reg_rva_out_Push_mioi_iswt0_cse <= and_572_cse;
      reg_start_PopNB_mioi_iswt0_cse <= and_574_rmff;
      reg_act_port_Push_mioi_iswt0_cse <= and_576_cse;
      reg_rva_in_PopNB_mioi_iswt0_cse <= fsm_output;
      pe_config_manager_counter_sva_dfm_3_1 <= MUX_v_4_2_2(4'b0000, operator_4_false_acc_nl,
          pe_config_UpdateManagerCounter_if_not_7_nl);
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= ~((pe_config_input_counter_sva_mx1 != (operator_16_false_acc_sdt_sva_1[7:0]))
          | (operator_16_false_acc_sdt_sva_1[8]));
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
      while_stage_0_3 <= reg_rva_in_PopNB_mioi_iswt0_cse;
      while_stage_0_4 <= while_stage_0_3;
      while_stage_0_5 <= while_stage_0_4;
      while_stage_0_6 <= while_stage_0_5;
      while_stage_0_7 <= while_stage_0_6;
      while_stage_0_8 <= while_stage_0_7;
      while_stage_0_9 <= while_stage_0_8;
      while_stage_0_10 <= while_stage_0_9;
      while_stage_0_11 <= while_stage_0_10;
      while_stage_0_12 <= while_stage_0_11;
      while_stage_0_13 <= while_stage_0_12;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_359_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[2];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_153_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[1];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_141_itm_1 <= pe_manager_base_weight_sva_mx3_0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1 <= ~ (pe_manager_base_weight_sva_mx1_3_0[2]);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_5_itm_1 <= ~ pe_manager_base_weight_sva_mx3_0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_4_itm_1 <= ~ (pe_manager_base_weight_sva_mx1_3_0[1]);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_1
          <= ~((pe_manager_base_weight_sva_mx1_3_0[2:1]!=2'b00) | pe_manager_base_weight_sva_mx3_0);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1 <= (pe_manager_base_weight_sva_mx1_3_0[2:1]==2'b11)
          & pe_manager_base_weight_sva_mx3_0 & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 <= (pe_manager_base_weight_sva_mx1_3_0[2:1]==2'b11)
          & (~ pe_manager_base_weight_sva_mx3_0) & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_1 <= (pe_manager_base_weight_sva_mx1_3_0[2])
          & pe_manager_base_weight_sva_mx3_0 & (~ (pe_manager_base_weight_sva_mx1_3_0[1]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      input_read_addrs_sva_1_1 <= nl_input_read_addrs_sva_1_1[7:0];
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
      weight_port_read_out_data_0_1_sva_15 <= weight_port_read_out_data_0_1_sva_mx0_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_11 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_11 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_11 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_2_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_10 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_11 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_11 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_11 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_11 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_191_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_11 <= rva_out_reg_data_15_9_sva_dfm_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_9 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_192_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_9 <= rva_out_reg_data_23_17_sva_dfm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_255_240_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_193_enex5 ) begin
      rva_out_reg_data_255_240_sva_dfm_4_6 <= rva_out_reg_data_255_240_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_239_224_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_194_enex5 ) begin
      rva_out_reg_data_239_224_sva_dfm_4_6 <= rva_out_reg_data_239_224_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_223_208_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_195_enex5 ) begin
      rva_out_reg_data_223_208_sva_dfm_4_6 <= rva_out_reg_data_223_208_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_207_192_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_196_enex5 ) begin
      rva_out_reg_data_207_192_sva_dfm_4_6 <= rva_out_reg_data_207_192_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_191_176_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_197_enex5 ) begin
      rva_out_reg_data_191_176_sva_dfm_4_6 <= rva_out_reg_data_191_176_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_175_160_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_198_enex5 ) begin
      rva_out_reg_data_175_160_sva_dfm_4_6 <= rva_out_reg_data_175_160_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_159_144_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_199_enex5 ) begin
      rva_out_reg_data_159_144_sva_dfm_4_6 <= rva_out_reg_data_159_144_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_143_128_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_200_enex5 ) begin
      rva_out_reg_data_143_128_sva_dfm_4_6 <= rva_out_reg_data_143_128_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_201_enex5 ) begin
      rva_out_reg_data_127_112_sva_dfm_4_6 <= rva_out_reg_data_127_112_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_96_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_202_enex5 ) begin
      rva_out_reg_data_111_96_sva_dfm_4_6 <= rva_out_reg_data_111_96_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_80_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_203_enex5 ) begin
      rva_out_reg_data_95_80_sva_dfm_4_6 <= rva_out_reg_data_95_80_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_6 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_204_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_6 <= rva_out_reg_data_39_36_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_4_6 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_205_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_4_6 <= rva_out_reg_data_79_64_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_6 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_206_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_6 <= rva_out_reg_data_46_40_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_63_sva_dfm_4_6 <= 1'b0;
      rva_out_reg_data_47_sva_dfm_4_6 <= 1'b0;
      input_read_req_valid_lpi_1_dfm_1_11 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9 <= 1'b0;
      rva_out_reg_data_35_32_sva_dfm_4_6_rsp_0 <= 2'b00;
      rva_out_reg_data_35_32_sva_dfm_4_6_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_29_cse ) begin
      rva_out_reg_data_63_sva_dfm_4_6 <= rva_out_reg_data_63_sva_dfm_4_5;
      rva_out_reg_data_47_sva_dfm_4_6 <= rva_out_reg_data_47_sva_dfm_4_5;
      input_read_req_valid_lpi_1_dfm_1_11 <= input_read_req_valid_lpi_1_dfm_1_10;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_9 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8;
      rva_out_reg_data_35_32_sva_dfm_4_6_rsp_0 <= rva_out_reg_data_35_32_sva_dfm_4_5_3_2;
      rva_out_reg_data_35_32_sva_dfm_4_6_rsp_1 <= rva_out_reg_data_35_32_sva_dfm_4_5_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_4_6 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_207_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_4_6 <= rva_out_reg_data_62_48_sva_dfm_4_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_6 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_6 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_6
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_6
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_6
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_6 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_6 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_6
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_6
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_6
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_6 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_172_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_6 <= weight_port_read_out_data_0_0_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_7_1_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_15_9_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_23_17_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_30_25_sva_dfm_6_5_2_1 <= 4'b0000;
      rva_out_reg_data_30_25_sva_dfm_6_1_0_1 <= 2'b00;
      rva_out_reg_data_0_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_8_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_16_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_31_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_24_sva_dfm_6 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_cse ) begin
      rva_out_reg_data_7_1_sva_dfm_6 <= rva_out_reg_data_7_1_sva_dfm_7;
      rva_out_reg_data_15_9_sva_dfm_6 <= rva_out_reg_data_15_9_sva_dfm_7;
      rva_out_reg_data_23_17_sva_dfm_6 <= rva_out_reg_data_23_17_sva_dfm_7;
      rva_out_reg_data_30_25_sva_dfm_6_5_2_1 <= rva_out_reg_data_30_25_sva_dfm_7_5_2;
      rva_out_reg_data_30_25_sva_dfm_6_1_0_1 <= rva_out_reg_data_30_25_sva_dfm_7_1_0;
      rva_out_reg_data_0_sva_dfm_6 <= rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_0_mx0;
      rva_out_reg_data_8_sva_dfm_6 <= rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_8_mx0;
      rva_out_reg_data_16_sva_dfm_6 <= rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_16_mx0;
      rva_out_reg_data_31_sva_dfm_6 <= rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_31_mx0;
      rva_out_reg_data_24_sva_dfm_6 <= rva_out_Push_mioi_m_data_rsc_dat_PECoreRun_24_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_6
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_57_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_6
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_6
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_58_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_6
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_125_cse ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd <= weight_port_read_out_data_0_1_sva_dfm_5_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_173_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_6_ftd_1 <= weight_port_read_out_data_0_1_sva_dfm_5_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_6
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_59_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_6
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_6
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_60_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_6
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_11 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11
          <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_cse ) begin
      rva_in_reg_rw_sva_11 <= rva_in_reg_rw_sva_10;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_11
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_11 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_6 ) begin
      rva_in_reg_rw_sva_st_1_11 <= rva_in_reg_rw_sva_st_1_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_11
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_11
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_9
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_11
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_11
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_255_224_sva_dfm_1_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_24 & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10
        ) begin
      act_port_reg_data_255_224_sva_dfm_1_1 <= act_port_reg_data_255_224_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_11 <= 1'b0;
      PECore_RunMac_PECore_RunMac_if_and_svs_11 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_11 <= 1'b0;
    end
    else if ( PECore_PushOutput_if_and_cse ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_11 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10;
      PECore_RunMac_PECore_RunMac_if_and_svs_11 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_10;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_11 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_31_0_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_63_32_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_95_64_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_127_96_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_159_128_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_191_160_sva <= 32'b00000000000000000000000000000000;
      act_port_reg_data_223_192_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( and_1072_cse ) begin
      act_port_reg_data_31_0_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_31_0_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_25_nl);
      act_port_reg_data_63_32_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_63_32_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_26_nl);
      act_port_reg_data_95_64_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_95_64_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_27_nl);
      act_port_reg_data_127_96_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_127_96_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_28_nl);
      act_port_reg_data_159_128_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_159_128_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_29_nl);
      act_port_reg_data_191_160_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_191_160_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_30_nl);
      act_port_reg_data_223_192_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_223_192_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_19_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_11 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_24 & (PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10
        | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10)) ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_11 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_10;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_6_35_0_sva <= 36'b000000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_24_enex5 ) begin
      accum_vector_data_6_35_0_sva <= accum_vector_data_6_35_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_5_35_0_sva <= 36'b000000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_25_enex5 ) begin
      accum_vector_data_5_35_0_sva <= accum_vector_data_5_35_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_4_35_0_sva <= 36'b000000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_26_enex5 ) begin
      accum_vector_data_4_35_0_sva <= accum_vector_data_4_35_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_3_35_0_sva <= 36'b000000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_27_enex5 ) begin
      accum_vector_data_3_35_0_sva <= accum_vector_data_3_35_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_2_35_0_sva <= 36'b000000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_28_enex5 ) begin
      accum_vector_data_2_35_0_sva <= accum_vector_data_2_35_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_1_35_0_sva <= 36'b000000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_29_enex5 ) begin
      accum_vector_data_1_35_0_sva <= accum_vector_data_1_35_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_0_35_0_sva <= 36'b000000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_30_enex5 ) begin
      accum_vector_data_0_35_0_sva <= accum_vector_data_0_35_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_10 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9
        | PECore_RunMac_PECore_RunMac_if_and_svs_st_9)) & while_stage_0_11 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_10 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_10 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_10 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_10 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_1_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_10 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_9;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_10 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_9;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_10 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_6_35_0_sva_dfm_1_1 <= 36'b000000000000000000000000000000000000;
      accum_vector_data_5_35_0_sva_dfm_1_1 <= 36'b000000000000000000000000000000000000;
      accum_vector_data_4_35_0_sva_dfm_1_1 <= 36'b000000000000000000000000000000000000;
      accum_vector_data_3_35_0_sva_dfm_1_1 <= 36'b000000000000000000000000000000000000;
      accum_vector_data_2_35_0_sva_dfm_1_1 <= 36'b000000000000000000000000000000000000;
      accum_vector_data_1_35_0_sva_dfm_1_1 <= 36'b000000000000000000000000000000000000;
      accum_vector_data_0_35_0_sva_dfm_1_1 <= 36'b000000000000000000000000000000000000;
    end
    else if ( and_1099_cse ) begin
      accum_vector_data_6_35_0_sva_dfm_1_1 <= MUX_v_36_2_2(36'b000000000000000000000000000000000000,
          PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_nl, PECore_UpdateFSM_switch_lp_not_31_nl);
      accum_vector_data_5_35_0_sva_dfm_1_1 <= MUX_v_36_2_2(36'b000000000000000000000000000000000000,
          PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_1_nl, PECore_UpdateFSM_switch_lp_not_32_nl);
      accum_vector_data_4_35_0_sva_dfm_1_1 <= MUX_v_36_2_2(36'b000000000000000000000000000000000000,
          PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_2_nl, PECore_UpdateFSM_switch_lp_not_33_nl);
      accum_vector_data_3_35_0_sva_dfm_1_1 <= MUX_v_36_2_2(36'b000000000000000000000000000000000000,
          PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_3_nl, PECore_UpdateFSM_switch_lp_not_34_nl);
      accum_vector_data_2_35_0_sva_dfm_1_1 <= MUX_v_36_2_2(36'b000000000000000000000000000000000000,
          PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_4_nl, PECore_UpdateFSM_switch_lp_not_35_nl);
      accum_vector_data_1_35_0_sva_dfm_1_1 <= MUX_v_36_2_2(36'b000000000000000000000000000000000000,
          PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_5_nl, PECore_UpdateFSM_switch_lp_not_36_nl);
      accum_vector_data_0_35_0_sva_dfm_1_1 <= MUX_v_36_2_2(36'b000000000000000000000000000000000000,
          PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_6_nl, PECore_UpdateFSM_switch_lp_not_21_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_10
          <= 1'b0;
      rva_in_reg_rw_sva_10 <= 1'b0;
    end
    else if ( while_if_and_6_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_10
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9;
      rva_in_reg_rw_sva_10 <= rva_in_reg_rw_sva_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_35_0_sva <= 36'b000000000000000000000000000000000000;
    end
    else if ( accum_vector_data_and_7_enex5 ) begin
      accum_vector_data_7_35_0_sva <= accum_vector_data_7_35_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
        | PECore_RunMac_PECore_RunMac_if_and_svs_st_8)) & while_stage_0_10 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_9 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_9 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_2_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_9 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_35_0_sva_dfm_1_1 <= 36'b000000000000000000000000000000000000;
    end
    else if ( and_1120_tmp ) begin
      accum_vector_data_7_35_0_sva_dfm_1_1 <= MUX_v_36_2_2(36'b000000000000000000000000000000000000,
          PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_7_nl, PECore_UpdateFSM_switch_lp_not_10_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9
          <= 1'b0;
      rva_in_reg_rw_sva_9 <= 1'b0;
    end
    else if ( while_if_and_7_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_9
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
      rva_in_reg_rw_sva_9 <= rva_in_reg_rw_sva_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
        | PECore_RunMac_PECore_RunMac_if_and_svs_st_7)) & while_stage_0_9 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_3_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= 1'b0;
      rva_in_reg_rw_sva_8 <= 1'b0;
    end
    else if ( while_if_and_8_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
      rva_in_reg_rw_sva_8 <= rva_in_reg_rw_sva_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_4_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= 1'b0;
      weight_port_read_out_data_0_3_sva <= 16'b0000000000000000;
      weight_port_read_out_data_0_2_sva <= 16'b0000000000000000;
      rva_in_reg_rw_sva_7 <= 1'b0;
      weight_port_read_out_data_0_1_sva_14_0 <= 15'b000000000000000;
    end
    else if ( while_if_and_9_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
      weight_port_read_out_data_0_3_sva <= weight_port_read_out_data_0_3_sva_mx0;
      weight_port_read_out_data_0_2_sva <= weight_port_read_out_data_0_2_sva_mx0;
      rva_in_reg_rw_sva_7 <= rva_in_reg_rw_sva_6;
      weight_port_read_out_data_0_1_sva_14_0 <= weight_port_read_out_data_0_1_sva_mx0_14_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_127_tmp ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_0_sva_dfm_1_mx0w0,
          weight_port_read_out_data_0_0_sva_dfm_mx0w1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1 <= 16'b0000000000000000;
    end
    else if ( mux_354_nl & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_0_2_sva_dfm_1_1 <= MUX1HOT_v_16_9_2(weight_port_read_out_data_0_2_sva_mx0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[31:16]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
          , weight_mem_run_3_for_5_and_166_nl , weight_mem_run_3_for_5_and_167_nl
          , weight_mem_run_3_for_5_and_168_nl , weight_mem_run_3_for_5_and_169_nl
          , weight_mem_run_3_for_5_and_170_nl , weight_mem_run_3_for_5_and_163_cse
          , weight_mem_run_3_for_5_and_172_nl});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1 <= 16'b0000000000000000;
    end
    else if ( mux_355_nl & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_1 <= MUX1HOT_v_16_9_2(weight_port_read_out_data_0_3_sva_mx0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[47:32]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
          , weight_mem_run_3_for_5_and_174_nl , weight_mem_run_3_for_5_and_175_nl
          , weight_mem_run_3_for_5_and_176_nl , weight_mem_run_3_for_5_and_177_nl
          , weight_mem_run_3_for_5_and_162_cse , weight_mem_run_3_for_5_and_179_nl
          , weight_mem_run_3_for_5_and_180_nl});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_5_mux_4_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_5_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_6_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_7_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_8_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_9_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_12_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_13_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_14_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_15_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_96_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_97_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_98_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_99_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_110_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_111_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_16_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_17_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_18_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_19_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_20_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_21_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_22_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_23_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_24_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_25_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_26_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_27_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_28_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_29_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_30_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_80_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_81_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_82_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_83_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_84_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_85_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_86_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_87_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_88_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_89_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_90_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_91_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_92_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_93_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_47_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_79_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_48_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_49_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_50_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_51_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_52_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_53_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_54_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_55_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_56_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_57_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_58_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_59_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_60_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_61_itm_1 <= 16'b0000000000000000;
      weight_mem_run_3_for_5_mux_62_itm_1 <= 16'b0000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_cse ) begin
      weight_mem_run_3_for_5_mux_4_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_4_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_5_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_5_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_6_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_6_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_7_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_7_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_8_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_8_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_9_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_9_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_12_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_12_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_13_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_13_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_14_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_14_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_15_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_0_15_sva_dfm_2,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011,
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_96_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_97_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_1_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_98_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_99_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_110_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_14_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_111_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_6_15_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_16_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_17_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_1_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_18_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_19_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_20_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_21_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_22_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_23_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_24_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_8_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_25_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_9_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_26_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_10_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_27_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_11_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_28_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_12_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_29_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_13_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_30_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_1_14_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_80_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_81_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_1_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_82_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_83_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_84_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_85_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_86_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_87_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_88_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_8_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_89_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_9_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_90_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_10_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_91_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_11_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_92_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_12_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_93_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_5_13_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013,
          weight_mem_run_3_for_land_6_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_47_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_2_15_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_mem_run_3_for_land_3_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_79_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_4_15_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_48_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_0_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_49_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_1_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_50_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_51_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_52_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_53_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_54_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_55_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_56_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_8_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_57_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_9_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_58_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_10_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_59_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_11_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_60_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_12_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_61_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_13_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_62_itm_1 <= MUX_v_16_2_2(weight_port_read_out_data_3_14_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_15_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_enex5 ) begin
      weight_port_read_out_data_1_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
          <= 16'b0000000000000000;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
          <= MUX_v_16_2_2(16'b0000000000000000, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_2_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_3 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= 1'b0;
      rva_in_reg_rw_sva_6 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_cse ) begin
      weight_mem_run_3_for_land_2_lpi_1_dfm_3 <= weight_mem_run_3_for_land_2_lpi_1_dfm_2;
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= weight_mem_run_3_for_land_3_lpi_1_dfm_2;
      weight_mem_run_3_for_land_5_lpi_1_dfm_3 <= weight_mem_run_3_for_land_5_lpi_1_dfm_2;
      weight_mem_run_3_for_land_4_lpi_1_dfm_3 <= weight_mem_run_3_for_land_4_lpi_1_dfm_2;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
      rva_in_reg_rw_sva_6 <= rva_in_reg_rw_sva_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_174_enex5 ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014
          <= 16'b0000000000000000;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[15:0]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[31:16]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[47:32]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[63:48]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[79:64]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[95:80]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[111:96]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[143:128]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[143:128]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[143:128]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[143:128]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[127:112]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[159:144]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[159:144]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[159:144]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[159:144]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[143:128]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[175:160]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[175:160]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[175:160]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[175:160]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[159:144]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[191:176]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[191:176]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[191:176]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[191:176]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[175:160]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[207:192]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[207:192]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[207:192]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[207:192]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[191:176]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[223:208]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[223:208]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[223:208]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[223:208]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[207:192]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[239:224]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[239:224]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[239:224]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[239:224]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[223:208]), {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_175_enex5 ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_176_enex5 ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_3_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_177_enex5 ) begin
      weight_port_read_out_data_2_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_4_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_178_enex5 ) begin
      weight_port_read_out_data_2_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_5_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_179_enex5 ) begin
      weight_port_read_out_data_2_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_6_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_180_enex5 ) begin
      weight_port_read_out_data_2_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_7_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_181_enex5 ) begin
      weight_port_read_out_data_2_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_8_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_182_enex5 ) begin
      weight_port_read_out_data_2_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_9_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_183_enex5 ) begin
      weight_port_read_out_data_2_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_10_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_184_enex5 ) begin
      weight_port_read_out_data_2_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_11_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_185_enex5 ) begin
      weight_port_read_out_data_2_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_12_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_186_enex5 ) begin
      weight_port_read_out_data_2_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_13_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_187_enex5 ) begin
      weight_port_read_out_data_2_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_14_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_188_enex5 ) begin
      weight_port_read_out_data_2_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_189_enex5 ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012
          <= 16'b0000000000000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014
          <= 16'b0000000000000000;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:0]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:0]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:0]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
          {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:16]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:16]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:16]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:16]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[15:0]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:32]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:32]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:32]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:32]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[31:16]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:48]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:48]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:48]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:48]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[47:32]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[79:64]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[79:64]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[79:64]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[79:64]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[79:64]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[63:48]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[95:80]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[95:80]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[95:80]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[95:80]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[95:80]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[79:64]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[111:96]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[111:96]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[111:96]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[111:96]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[111:96]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[95:80]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[127:112]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[127:112]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[127:112]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[127:112]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[127:112]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[111:96]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[143:128]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[143:128]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[143:128]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[143:128]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[143:128]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[127:112]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[159:144]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[159:144]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[159:144]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[159:144]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[159:144]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[143:128]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[175:160]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[175:160]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[175:160]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[175:160]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[175:160]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[159:144]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[191:176]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[191:176]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[191:176]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[191:176]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[191:176]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[175:160]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[207:192]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[207:192]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[207:192]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[207:192]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[207:192]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[191:176]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[223:208]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[223:208]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[223:208]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[223:208]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[223:208]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[207:192]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014
          <= MUX_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[239:224]),
          (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[239:224]),
          (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[239:224]),
          (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[239:224]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[239:224]),
          (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[223:208]), {weight_read_addrs_4_14_2_lpi_1_dfm_3_0
          , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_1_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_190_enex5 ) begin
      weight_port_read_out_data_4_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_2_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_191_enex5 ) begin
      weight_port_read_out_data_4_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_3_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_192_enex5 ) begin
      weight_port_read_out_data_4_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_4_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_193_enex5 ) begin
      weight_port_read_out_data_4_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_5_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_194_enex5 ) begin
      weight_port_read_out_data_4_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_6_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_195_enex5 ) begin
      weight_port_read_out_data_4_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_7_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_196_enex5 ) begin
      weight_port_read_out_data_4_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_8_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_197_enex5 ) begin
      weight_port_read_out_data_4_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_9_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_198_enex5 ) begin
      weight_port_read_out_data_4_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_10_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_199_enex5 ) begin
      weight_port_read_out_data_4_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_11_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_200_enex5 ) begin
      weight_port_read_out_data_4_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_12_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_201_enex5 ) begin
      weight_port_read_out_data_4_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_13_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_202_enex5 ) begin
      weight_port_read_out_data_4_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_14_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_203_enex5 ) begin
      weight_port_read_out_data_4_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_15_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_31_enex5 ) begin
      weight_port_read_out_data_3_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
          <= 16'b0000000000000000;
    end
    else if ( data_in_tmp_operator_2_for_and_31_tmp ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000
          <= MUX_v_16_2_2(16'b0000000000000000, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_1_nl,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_5_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_5,
          (weight_port_read_out_data_0_3_sva_dfm_2[15]), PECore_PushAxiRsp_if_else_mux_26_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_46_tmp , while_and_45_cse});
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5,
          (weight_port_read_out_data_0_2_sva_dfm_2[15]), PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_46_tmp , while_and_45_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_1)
        & while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1)
        & while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_5 <= 1'b0;
      rva_in_reg_rw_sva_st_5 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_2_cse ) begin
      rva_in_reg_rw_sva_st_1_5 <= rva_in_reg_rw_sva_st_1_4;
      rva_in_reg_rw_sva_st_5 <= rva_in_reg_rw_sva_st_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_1_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2 <= 1'b0;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= 1'b0;
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_run_3_for_5_and_140_itm_2 <= 1'b0;
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_run_3_for_5_and_142_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_143_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_144_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_132_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_135_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_126_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1 <= 1'b0;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= 3'b000;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_12_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_14_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_15_itm_1_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_16_itm_1_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_6_itm_1_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_7_itm_2_cse <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_2 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_146_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_147_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_148_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_149_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_151_itm_2 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_152_itm_2_cse <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_6_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= MUX_v_256_2_2(weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= MUX_v_256_2_2(weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= MUX_v_256_2_2(weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_run_3_for_5_and_140_itm_2 <= weight_mem_run_3_for_5_and_140_itm_1;
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= MUX_v_256_2_2(weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_run_3_for_5_and_142_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_143_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_144_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b111)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_132_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b011)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_135_itm_2 <= weight_mem_run_3_for_5_and_135_itm_1;
      weight_mem_run_3_for_5_and_126_itm_2 <= weight_mem_run_3_for_5_and_126_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_2_2_0!=3'b000));
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= weight_read_addrs_7_lpi_1_dfm_2_2_0;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
      reg_weight_mem_run_3_for_5_and_12_itm_2_cse <= weight_mem_run_3_for_5_and_12_itm_1;
      reg_weight_mem_run_3_for_5_and_14_itm_2_cse <= weight_mem_run_3_for_5_and_14_itm_1;
      reg_weight_mem_run_3_for_5_and_15_itm_1_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1;
      reg_weight_mem_run_3_for_5_and_16_itm_1_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1_1;
      reg_weight_mem_run_3_for_5_and_6_itm_1_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_278_itm_1;
      reg_weight_mem_run_3_for_5_and_7_itm_2_cse <= weight_mem_run_3_for_5_and_7_itm_1;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= weight_read_addrs_5_lpi_1_dfm_2_2_0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1;
      reg_weight_mem_run_3_for_5_and_146_itm_2_cse <= weight_mem_run_3_for_5_and_146_itm_1;
      reg_weight_mem_run_3_for_5_and_147_itm_2_cse <= weight_mem_run_3_for_5_and_147_itm_1;
      reg_weight_mem_run_3_for_5_and_148_itm_2_cse <= weight_mem_run_3_for_5_and_148_itm_1;
      reg_weight_mem_run_3_for_5_and_149_itm_2_cse <= weight_mem_run_3_for_5_and_149_itm_1;
      weight_mem_run_3_for_5_and_150_itm_2 <= weight_mem_run_3_for_5_and_150_itm_1;
      weight_mem_run_3_for_5_and_151_itm_2 <= weight_mem_run_3_for_5_and_151_itm_1;
      reg_weight_mem_run_3_for_5_and_152_itm_2_cse <= weight_mem_run_3_for_5_and_152_itm_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_15_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1130_cse | or_dcpl_753 | or_dcpl_752) & and_dcpl_808 & PECoreRun_wen
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_15_sva_dfm_1 <= weight_port_read_out_data_7_15_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_14_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1135_cse | weight_mem_run_3_for_5_and_135_itm_2 | weight_mem_run_3_for_5_and_142_itm_1
        | weight_mem_run_3_for_5_and_132_itm_1) & and_dcpl_808 & PECoreRun_wen &
        (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_14_sva_dfm_1 <= weight_port_read_out_data_7_14_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_13_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_7_11_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_7_7_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( and_1141_cse ) begin
      weight_port_read_out_data_7_13_sva_dfm_1 <= weight_port_read_out_data_7_13_sva_dfm_3;
      weight_port_read_out_data_7_11_sva_dfm_1 <= weight_port_read_out_data_7_11_sva_dfm_3;
      weight_port_read_out_data_7_7_sva_dfm_1 <= weight_port_read_out_data_7_7_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_12_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1130_cse | or_dcpl_766 | weight_mem_run_3_for_5_and_142_itm_1
        | weight_mem_run_3_for_5_and_132_itm_1) & and_dcpl_808 & PECoreRun_wen &
        (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_12_sva_dfm_1 <= weight_port_read_out_data_7_12_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_10_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_7_9_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( and_1156_cse ) begin
      weight_port_read_out_data_7_10_sva_dfm_1 <= weight_port_read_out_data_7_10_sva_dfm_3;
      weight_port_read_out_data_7_9_sva_dfm_1 <= weight_port_read_out_data_7_9_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_8_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1165_cse | weight_mem_run_3_for_5_and_143_itm_1 | weight_mem_run_3_for_5_and_142_itm_1
        | weight_mem_run_3_for_5_and_140_itm_2) & and_dcpl_808 & PECoreRun_wen &
        (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_8_sva_dfm_1 <= weight_port_read_out_data_7_8_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_6_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1135_cse | or_dcpl_792 | weight_mem_run_3_for_5_and_140_itm_2)
        & and_dcpl_808 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_6_sva_dfm_1 <= weight_port_read_out_data_7_6_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_5_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1130_cse | or_dcpl_766 | or_dcpl_752) & and_dcpl_808 & PECoreRun_wen
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_5_sva_dfm_1 <= weight_port_read_out_data_7_5_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_4_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1165_cse | or_dcpl_792 | weight_mem_run_3_for_5_and_132_itm_1)
        & and_dcpl_808 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_4_sva_dfm_1 <= weight_port_read_out_data_7_4_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_3_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1165_cse | or_dcpl_761 | weight_mem_run_3_for_5_and_132_itm_1)
        & and_dcpl_808 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_3_sva_dfm_1 <= weight_port_read_out_data_7_3_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_2_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1130_cse | or_dcpl_766 | weight_mem_run_3_for_5_and_126_itm_2
        | weight_mem_run_3_for_5_and_132_itm_1) & and_dcpl_808 & PECoreRun_wen &
        (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_7_2_sva_dfm_1 <= weight_port_read_out_data_7_2_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_1_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_7_0_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( and_1201_cse ) begin
      weight_port_read_out_data_7_1_sva_dfm_1 <= weight_port_read_out_data_7_1_sva_dfm_3;
      weight_port_read_out_data_7_0_sva_dfm_1 <= weight_port_read_out_data_7_0_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= 1'b0;
      rva_in_reg_rw_sva_5 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_5_cse ) begin
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= weight_mem_run_3_for_land_1_lpi_1_dfm_2;
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= weight_mem_run_3_for_land_7_lpi_1_dfm_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= weight_mem_run_3_for_land_3_lpi_1_dfm_1;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= weight_mem_run_3_for_land_5_lpi_1_dfm_1;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
      rva_in_reg_rw_sva_5 <= rva_in_reg_rw_sva_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_15_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1210_cse | reg_weight_mem_run_3_for_5_and_16_itm_1_cse | reg_weight_mem_run_3_for_5_and_15_itm_1_cse
        | reg_weight_mem_run_3_for_5_and_14_itm_2_cse | reg_weight_mem_run_3_for_5_and_12_itm_2_cse)
        & and_dcpl_808 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_5_15_sva_dfm_1 <= weight_port_read_out_data_5_15_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_14_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (and_1210_cse | reg_weight_mem_run_3_for_5_and_16_itm_1_cse | reg_weight_mem_run_3_for_5_and_7_itm_2_cse
        | reg_weight_mem_run_3_for_5_and_6_itm_1_cse | reg_weight_mem_run_3_for_5_and_12_itm_2_cse)
        & and_dcpl_808 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_5_14_sva_dfm_1 <= weight_port_read_out_data_5_14_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= 16'b0000000000000000;
    end
    else if ( mux_376_nl & and_dcpl_808 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & mux_5_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1
          <= MUX_v_16_2_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[15:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_48_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & mux_6_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_256U_2_for_1_marshaller_AddField_ac_int_16_false_16_11_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_15_0_1_itm_1
          <= MUX_v_16_2_2((weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[15:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_80_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_255_16 <= 240'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_633 | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & ((~(while_stage_0_6 & weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_255_16 <= weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[255:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_633 | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & ((~(while_stage_0_6 & weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_RunFSM_switch_lp_equal_tmp_1_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_UpdateFSM_switch_lp_equal_tmp_2_3 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_empty_sva_1[2])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_7_nl) & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_380_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_2_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_76 & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]))
        ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_76 & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= 1'b0;
      rva_in_reg_rw_sva_4 <= 1'b0;
    end
    else if ( while_if_and_12_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_125_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3_1
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3_1
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1_1
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1_1);
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp |
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp |
          Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3_1);
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & weight_mem_read_arbxbar_xbar_1_for_3_8_for_7_or_cse;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
      rva_in_reg_rw_sva_4 <= rva_in_reg_rw_sva_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_52_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_58_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse & (and_dcpl_76 | Arbiter_8U_Roundrobin_pick_and_14_cse)
        & or_dcpl_47 ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0,
          Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1, Arbiter_8U_Roundrobin_pick_and_14_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_64_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse & (and_dcpl_76 | Arbiter_8U_Roundrobin_pick_and_13_cse)
        & or_dcpl_48 ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0,
          Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1, Arbiter_8U_Roundrobin_pick_and_13_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_69_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse & (and_dcpl_76 | Arbiter_8U_Roundrobin_pick_and_44_cse)
        & or_dcpl_50 ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_80_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1, Arbiter_8U_Roundrobin_pick_and_44_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_74_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_79_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse & (and_dcpl_76 | Arbiter_8U_Roundrobin_pick_and_8_cse)
        & or_dcpl_53 ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0,
          Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1, Arbiter_8U_Roundrobin_pick_and_8_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_85_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_90_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= weight_mem_read_arbxbar_arbiters_next_0_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva <= 15'b000000000000000;
    end
    else if ( (~ mux_378_nl) & fsm_output & while_stage_0_5 & PECoreRun_wen ) begin
      pe_manager_base_weight_sva <= pe_manager_base_weight_sva_mx2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= 11'b00000000000;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= 1'b0;
    end
    else if ( weight_read_addrs_and_4_cse ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= MUX_v_11_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl,
          weight_read_addrs_0_14_4_lpi_1_dfm_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= MUX_s_1_2_2((weight_read_addrs_0_3_0_lpi_1_dfm_4[3]),
          (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]))) & while_stage_0_4 )
        begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= MUX_s_1_2_2((~ (pe_manager_base_weight_sva_mx1_3_0[1])), (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_48_enex5 ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_15_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_49_enex5 ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_14_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_50_enex5 ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_13_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_51_enex5 ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_12_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_52_enex5 ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_11_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_53_enex5 ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_10_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_54_enex5 ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_9_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_55_enex5 ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_8_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_56_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_57_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_58_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_59_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_60_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_61_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_62_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_63_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= 12'b000000000000;
    end
    else if ( weight_write_addrs_and_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= weight_write_addrs_lpi_1_dfm_1_2[14:3];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_133 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_133 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= 1'b0;
      weight_read_addrs_1_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_3_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= 13'b0000000000000;
      weight_read_addrs_5_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_7_lpi_1_dfm_1 <= 15'b000000000000000;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1,
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
      weight_read_addrs_1_lpi_1_dfm_1 <= weight_read_addrs_1_lpi_1_dfm_1_1;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_3_lpi_1_dfm_1 <= weight_read_addrs_3_lpi_1_dfm_1_1;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_1 <= weight_read_addrs_5_lpi_1_dfm_1_1;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_7_lpi_1_dfm_1 <= weight_read_addrs_7_lpi_1_dfm_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_5_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_5_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= or_185_cse;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
          & or_185_cse;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= Arbiter_8U_Roundrobin_pick_1_if_1_and_30_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_not_185,
          weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0, and_dcpl_588);
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0, and_115_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0,
          (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_5_tmp);
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0, and_122_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0,
          (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp);
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0,
          (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp);
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0,
          (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          or_185_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0,
          (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_363_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= 1'b0;
      rva_in_reg_rw_sva_3 <= 1'b0;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1 <= MUX_s_1_2_2((pe_manager_base_weight_sva_mx1_3_0[2]),
          reg_rva_in_reg_rw_sva_2_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_363_itm_1 <= MUX_s_1_2_2(pe_manager_base_weight_sva_mx3_0,
          reg_rva_in_reg_rw_sva_2_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      rva_in_reg_rw_sva_3 <= reg_rva_in_reg_rw_sva_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_31_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= 1'b0;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= 8'b00000000;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_1_for_and_cse ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_31_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b101)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b110)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= weight_mem_write_arbxbar_xbar_for_lshift_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_and_85_cse ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_590);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_590);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_590);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_590);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_590);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_590);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_590);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_590);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_64_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse & ((~ while_stage_0_5) | while_and_1282_itm_1)
        ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= MUX_v_15_2_2(pe_manager_base_weight_sva_mx2,
          PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1, while_and_1282_itm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_64_enex5 ) begin
      weight_write_data_data_0_15_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_15_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_65_enex5 ) begin
      weight_write_data_data_0_14_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_14_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_66_enex5 ) begin
      weight_write_data_data_0_13_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_13_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_67_enex5 ) begin
      weight_write_data_data_0_12_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_12_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_68_enex5 ) begin
      weight_write_data_data_0_11_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_11_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_69_enex5 ) begin
      weight_write_data_data_0_10_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_10_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_70_enex5 ) begin
      weight_write_data_data_0_9_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_9_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_71_enex5 ) begin
      weight_write_data_data_0_8_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_8_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_72_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_7_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_73_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_6_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_74_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_5_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_75_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_76_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_3_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_77_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_2_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_78_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_1_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= 16'b0000000000000000;
    end
    else if ( weight_write_data_data_and_79_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= 15'b000000000000000;
    end
    else if ( weight_write_addrs_and_3_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= weight_write_addrs_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( weight_write_data_data_and_16_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_2_cse <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= 1'b0;
      while_and_1282_itm_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_3_cse ) begin
      reg_rva_in_reg_rw_sva_2_cse <= reg_rva_in_reg_rw_sva_st_1_1_cse;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= MUX_s_1_2_2(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
      while_and_1282_itm_1 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1
          & PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
          & reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= 4'b0000;
    end
    else if ( weight_read_addrs_and_enex5 ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= 11'b00000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_176 ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_2_1_sva <= 2'b00;
      pe_config_is_zero_first_sva <= 1'b0;
    end
    else if ( state_and_cse ) begin
      state_2_1_sva <= state_mux_1_cse;
      pe_config_is_zero_first_sva <= pe_config_is_zero_first_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_0_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_637) ) begin
      state_0_sva <= PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_manager_counter_sva <= 4'b0000;
    end
    else if ( (((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:2]==6'b000000) & nor_518_cse
        & nor_520_cse & nor_521_cse & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])))
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & rva_in_PopNB_mioi_return_rsc_z_mxwt
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]==2'b00) & and_dcpl_183)
        | and_1227_cse) & PECoreRun_wen ) begin
      pe_config_manager_counter_sva <= MUX_v_4_2_2(pe_config_manager_counter_sva_dfm_3_1,
          PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl,
          and_622_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_num_manager_sva <= 4'b0001;
      pe_config_num_output_sva <= 8'b00000001;
    end
    else if ( pe_config_num_manager_and_cse ) begin
      pe_config_num_manager_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[35:32];
      pe_config_num_output_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= 1'b0;
      state_2_1_sva_dfm_1 <= 2'b00;
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= 8'b00000000;
      input_write_req_valid_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_4_cse ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= rva_in_PopNB_mioi_return_rsc_z_mxwt;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
      state_2_1_sva_dfm_1 <= MUX_v_2_2_2(PECore_UpdateFSM_switch_lp_and_1_nl, state_mux_1_cse,
          rva_in_PopNB_mioi_return_rsc_z_mxwt);
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= and_279_cse;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0];
      input_write_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= 1'b0;
      PECore_RunFSM_switch_lp_nor_tmp_1 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_9_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= PECore_UpdateFSM_switch_lp_equal_tmp_6;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= ~(PECore_RunScale_PECore_RunScale_if_and_1_svs_1
          | PECore_UpdateFSM_switch_lp_nor_tmp_1);
      PECore_RunFSM_switch_lp_nor_tmp_1 <= ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
          | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(or_142_cse | or_dcpl_637 | (~ fsm_output))) & (mux_115_cse
        | rva_in_PopNB_mioi_return_rsc_z_mxwt | (~ reg_rva_in_PopNB_mioi_iswt0_cse))
        ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= input_port_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva <= 8'b00000000;
    end
    else if ( or_1293_cse & mux_379_nl & weight_mem_read_arbxbar_arbiters_next_and_cse
        & while_stage_0_3 ) begin
      pe_config_input_counter_sva <= pe_config_input_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva <= 8'b00000000;
    end
    else if ( or_1293_cse & mux_380_nl & while_stage_0_3 & fsm_output & PECoreRun_wen
        ) begin
      pe_config_output_counter_sva <= pe_config_output_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      operator_8_false_acc_sdt_sva_1 <= 9'b000000000;
    end
    else if ( pe_config_UpdateManagerCounter_if_if_and_enex5 ) begin
      operator_8_false_acc_sdt_sva_1 <= nl_operator_8_false_acc_sdt_sva_1[8:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiWrite_switch_lp_and_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_255_224_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( mux_390_nl & fsm_output & while_stage_0_12 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_10)
        ) begin
      act_port_reg_data_255_224_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          act_port_reg_data_255_224_sva_dfm_3, PECore_UpdateFSM_switch_lp_not_11_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Datapath_for_6_ProductSum_for_acc_1_1 <= 34'b0000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
        & PECore_RunMac_PECore_RunMac_if_and_svs_st_8 & (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8)
        & while_stage_0_10 ) begin
      Datapath_for_6_ProductSum_for_acc_1_1 <= Datapath_for_4_ProductSum_for_acc_9_cmp_40_z;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_16_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_0_1_sva_dfm_1_14_0 <= 15'b000000000000000;
    end
    else if ( and_1266_cse ) begin
      weight_port_read_out_data_0_3_sva_dfm_1 <= weight_port_read_out_data_0_3_sva_dfm_2;
      weight_port_read_out_data_0_1_sva_dfm_1_14_0 <= MUX_v_15_2_2(15'b000000000000000,
          mux1h_7_nl, not_2496_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( (mux_396_nl | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_231_itm_1
        | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
        | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1) & and_dcpl_195
        & PECoreRun_wen ) begin
      weight_port_read_out_data_0_2_sva_dfm_1 <= weight_port_read_out_data_0_2_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & weight_mem_run_3_for_land_3_lpi_1_dfm_1 & while_stage_0_6
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= rva_out_reg_data_35_32_sva_dfm_1_4_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_36_nl & while_stage_0_6 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2 <= 2'b00;
    end
    else if ( weight_read_addrs_and_15_cse ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_itm_2 <= rva_out_reg_data_30_25_sva_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
      pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2 <= 1'b0;
    end
    else if ( weight_read_addrs_and_16_cse ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
      pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_2 <= pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_4_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_5_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_6_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_7_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_8_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_9_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_10_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_11_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_12_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_13_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_14_sva_dfm_2 <= 16'b0000000000000000;
      weight_port_read_out_data_0_15_sva_dfm_2 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_50_cse ) begin
      weight_port_read_out_data_0_4_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_63_48_sva_1,
          while_and_46_tmp);
      weight_port_read_out_data_0_5_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_79_64_sva_1,
          while_and_46_tmp);
      weight_port_read_out_data_0_6_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_95_80_sva_1,
          while_and_46_tmp);
      weight_port_read_out_data_0_7_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_111_9000000,
          while_and_46_tmp);
      weight_port_read_out_data_0_8_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_127_1000000,
          while_and_46_tmp);
      weight_port_read_out_data_0_9_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_143_1000000,
          while_and_46_tmp);
      weight_port_read_out_data_0_10_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_159_1000000,
          while_and_46_tmp);
      weight_port_read_out_data_0_11_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_175_1000000,
          while_and_46_tmp);
      weight_port_read_out_data_0_12_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_191_1000000,
          while_and_46_tmp);
      weight_port_read_out_data_0_13_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_207_1000000,
          while_and_46_tmp);
      weight_port_read_out_data_0_14_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_223_2000000,
          while_and_46_tmp);
      weight_port_read_out_data_0_15_sva_dfm_2 <= MUX_v_16_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_16_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_256_255_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_3_0_16_15_0_sdt_239_2000000,
          while_and_46_tmp);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_1_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_8_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_9_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_10_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_11_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_12_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_13_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_14_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_6_15_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_134_cse ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
      weight_port_read_out_data_6_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
      weight_port_read_out_data_6_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000;
      weight_port_read_out_data_6_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
      weight_port_read_out_data_6_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
      weight_port_read_out_data_6_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
      weight_port_read_out_data_6_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
      weight_port_read_out_data_6_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
      weight_port_read_out_data_6_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
      weight_port_read_out_data_6_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_1_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_2_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_3_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_4_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_5_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_6_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_7_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_8_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_9_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_10_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_11_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_12_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_13_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_1_14_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_78_cse ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
      weight_port_read_out_data_1_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
      weight_port_read_out_data_1_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
      weight_port_read_out_data_1_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
      weight_port_read_out_data_1_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
      weight_port_read_out_data_1_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
      weight_port_read_out_data_1_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
      weight_port_read_out_data_1_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
      weight_port_read_out_data_1_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
      weight_port_read_out_data_1_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
      weight_port_read_out_data_1_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
      weight_port_read_out_data_1_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
      weight_port_read_out_data_1_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
      weight_port_read_out_data_1_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
      weight_port_read_out_data_1_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_1_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_2_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_3_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_4_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_5_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_6_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_7_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_8_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_9_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_10_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_11_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_12_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_5_13_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_150_cse ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
      weight_port_read_out_data_5_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
      weight_port_read_out_data_5_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
      weight_port_read_out_data_5_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
      weight_port_read_out_data_5_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
      weight_port_read_out_data_5_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
      weight_port_read_out_data_5_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
      weight_port_read_out_data_5_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
      weight_port_read_out_data_5_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
      weight_port_read_out_data_5_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
      weight_port_read_out_data_5_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
      weight_port_read_out_data_5_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
      weight_port_read_out_data_5_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
      weight_port_read_out_data_5_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_6_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_15_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_run_3_for_land_3_lpi_1_dfm_2) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
        | (~ while_stage_0_7))) ) begin
      weight_port_read_out_data_2_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_15_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_633 | (~ weight_mem_run_3_for_land_5_lpi_1_dfm_2)
        | (~ fsm_output))) & ((~(while_stage_0_6 & weight_mem_run_3_for_land_5_lpi_1_dfm_1))
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        ) begin
      weight_port_read_out_data_4_15_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_0_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_1_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_2_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_3_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_4_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_5_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_6_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_7_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_8_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_9_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_10_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_11_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_12_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_13_sva_dfm_1 <= 16'b0000000000000000;
      weight_port_read_out_data_3_14_sva_dfm_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_109_cse ) begin
      weight_port_read_out_data_3_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000;
      weight_port_read_out_data_3_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000001;
      weight_port_read_out_data_3_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000002;
      weight_port_read_out_data_3_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000003;
      weight_port_read_out_data_3_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000004;
      weight_port_read_out_data_3_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000005;
      weight_port_read_out_data_3_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006;
      weight_port_read_out_data_3_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007;
      weight_port_read_out_data_3_8_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000008;
      weight_port_read_out_data_3_9_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000009;
      weight_port_read_out_data_3_10_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000010;
      weight_port_read_out_data_3_11_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000011;
      weight_port_read_out_data_3_12_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000012;
      weight_port_read_out_data_3_13_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000013;
      weight_port_read_out_data_3_14_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000014;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2 <= 16'b0000000000000000;
    end
    else if ( mux_399_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_0_sva_dfm_2 <= MUX_v_16_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w1,
          weight_port_read_out_data_0_0_sva_dfm_1_mx0w0, and_dcpl_45);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_336_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_328_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_336_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_328_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_37_nl & while_stage_0_6 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_36_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_374_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_36_itm_1
          <= ~((weight_read_addrs_5_lpi_1_dfm_2_2_0!=3'b000));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 <= 1'b0;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_378_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= weight_read_addrs_3_lpi_1_dfm_2_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_231_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_382_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_136_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_231_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_215_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_18_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_204_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_14_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_387_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_14_itm_1
          <= crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b110)
          & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1 <= 1'b0;
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_389_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_28_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_104_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_3
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_3 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_3 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_3 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_104_itm_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_100_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_3
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_5_and_140_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_135_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_126_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_14_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_12_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_7_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_152_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_151_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_149_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_148_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_147_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_146_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= 1'b0;
    end
    else if ( weight_read_addrs_and_19_cse ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= weight_read_addrs_7_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= weight_read_addrs_5_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_5_and_140_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_135_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_126_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_14_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1;
      weight_mem_run_3_for_5_and_12_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_weight_mem_run_3_for_and_5_tmp;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= ~((weight_read_addrs_5_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_7_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1;
      weight_mem_run_3_for_5_and_152_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1;
      weight_mem_run_3_for_5_and_151_itm_1 <= (pe_manager_base_weight_sva[2]) & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_380_itm_1
          & (~ (pe_manager_base_weight_sva[0])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_150_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1
          & (pe_manager_base_weight_sva[0]) & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_149_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
      weight_mem_run_3_for_5_and_148_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_40_itm_1;
      weight_mem_run_3_for_5_and_147_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
      weight_mem_run_3_for_5_and_146_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_18_itm_1 <= ~((pe_manager_base_weight_sva[2:1]!=2'b00)
          | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_363_itm_1);
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & ((~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        | (~ while_stage_0_6))) ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & ((~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_1284_cse | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
        | (~ fsm_output))) & ((~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_1284_cse | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
        | (~ fsm_output))) & mux_41_nl ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & ((~ weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_21_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_27_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= 1'b0;
    end
    else if ( operator_15_false_1_and_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        | (~ while_stage_0_4))) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~ or_185_cse) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        | (~ while_stage_0_4))) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(or_188_cse | (~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_2_tmp)))
        ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_3_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        | (~ while_stage_0_4))) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_122_cse | or_188_cse)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_5_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        | (~ while_stage_0_4))) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_115_cse | or_188_cse)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= 15'b000000000000000;
    end
    else if ( PEManager_15U_PEManagerWrite_and_enex5 ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= rva_in_reg_data_sva_1[30:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_num_input_sva <= 8'b00000001;
      pe_manager_base_bias_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_num_input_and_cse ) begin
      pe_manager_num_input_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      pe_manager_base_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[46:32];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_is_valid_sva <= 1'b0;
      pe_config_is_cluster_sva <= 1'b0;
      pe_config_is_bias_sva <= 1'b0;
    end
    else if ( pe_config_is_valid_and_cse ) begin
      pe_config_is_valid_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
      pe_config_is_cluster_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[16];
      pe_config_is_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_zero_active_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & and_279_cse & (~ PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)
        & (~ or_dcpl_648) ) begin
      pe_manager_zero_active_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva_dfm_1 <= 8'b00000000;
      pe_config_input_counter_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1294_cse ) begin
      pe_config_output_counter_sva_dfm_1 <= MUX_v_8_2_2(8'b00000000, pe_config_output_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
      pe_config_input_counter_sva_dfm_1 <= MUX_v_8_2_2(8'b00000000, pe_config_input_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_mux_27_itm_1 <= 1'b0;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= 4'b0000;
      weight_write_data_data_0_15_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_14_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_13_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_12_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_11_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_10_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_9_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_8_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= 16'b0000000000000000;
      weight_write_addrs_lpi_1_dfm_1_1 <= 15'b000000000000000;
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= 11'b00000000000;
    end
    else if ( while_if_and_16_cse ) begin
      while_if_mux_27_itm_1 <= MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_27_nl,
          rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:0])
          & ({{3{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_4_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
      weight_write_data_data_0_15_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[255:240])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_14_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[239:224])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_13_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[223:208])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_12_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[207:192])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_11_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[191:176])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_10_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[175:160])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_9_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[159:144])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_8_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[143:128])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:112])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:96])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:80])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:64])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:48])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:32])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:16])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:0])
          & ({{15{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{15{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_addrs_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:0])
          & ({{14{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{14{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:4])
          & ({{10{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_11_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
        | PECore_RunMac_PECore_RunMac_if_and_svs_st_6)) & while_stage_0_8 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_4 <= 1'b0;
      rva_in_reg_rw_sva_st_4 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_5_cse ) begin
      rva_in_reg_rw_sva_st_1_4 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_363_itm_1;
      rva_in_reg_rw_sva_st_4 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_376_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_10 <= 1'b0;
      rva_in_reg_rw_sva_st_10 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_6_cse ) begin
      rva_in_reg_rw_sva_st_1_10 <= rva_in_reg_rw_sva_st_1_9;
      rva_in_reg_rw_sva_st_10 <= rva_in_reg_rw_sva_st_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= 4'b0000;
    end
    else if ( PECoreRun_wen & and_dcpl_226 ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_9_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_5 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_5 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_61_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_62_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_63_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_64_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_2_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_10 <= 1'b0;
      rva_out_reg_data_47_sva_dfm_4_5 <= 1'b0;
      rva_out_reg_data_63_sva_dfm_4_5 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8 <= 1'b0;
      rva_out_reg_data_35_32_sva_dfm_4_5_3_2 <= 2'b00;
      rva_out_reg_data_35_32_sva_dfm_4_5_1_0 <= 2'b00;
    end
    else if ( input_read_req_valid_and_1_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_10 <= input_read_req_valid_lpi_1_dfm_1_9;
      rva_out_reg_data_47_sva_dfm_4_5 <= rva_out_reg_data_47_sva_dfm_4_4;
      rva_out_reg_data_63_sva_dfm_4_5 <= rva_out_reg_data_63_sva_dfm_4_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
      rva_out_reg_data_35_32_sva_dfm_4_5_3_2 <= reg_rva_out_reg_data_35_32_sva_dfm_4_4_ftd;
      rva_out_reg_data_35_32_sva_dfm_4_5_1_0 <= reg_rva_out_reg_data_35_32_sva_dfm_4_4_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_10 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_7_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_10 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_8_ftd <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_208_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_8_ftd <= rva_out_reg_data_30_25_sva_dfm_7_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_8_ftd_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_47_cse ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_8_ftd_1 <= rva_out_reg_data_30_25_sva_dfm_7_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_8 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_209_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_8 <= rva_out_reg_data_23_17_sva_dfm_7_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_10 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_210_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_10 <= rva_out_reg_data_15_9_sva_dfm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_5 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_204_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_5 <= weight_port_read_out_data_0_0_sva_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_5 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_211_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_5 <= rva_out_reg_data_39_36_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_212_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_5 <= rva_out_reg_data_46_40_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_4_5 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_213_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_4_5 <= rva_out_reg_data_62_48_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_255_240_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_214_enex5 ) begin
      rva_out_reg_data_255_240_sva_dfm_4_5 <= rva_out_reg_data_255_240_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_239_224_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_215_enex5 ) begin
      rva_out_reg_data_239_224_sva_dfm_4_5 <= rva_out_reg_data_239_224_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_223_208_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_216_enex5 ) begin
      rva_out_reg_data_223_208_sva_dfm_4_5 <= rva_out_reg_data_223_208_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_207_192_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_217_enex5 ) begin
      rva_out_reg_data_207_192_sva_dfm_4_5 <= rva_out_reg_data_207_192_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_191_176_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_218_enex5 ) begin
      rva_out_reg_data_191_176_sva_dfm_4_5 <= rva_out_reg_data_191_176_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_175_160_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_219_enex5 ) begin
      rva_out_reg_data_175_160_sva_dfm_4_5 <= rva_out_reg_data_175_160_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_159_144_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_220_enex5 ) begin
      rva_out_reg_data_159_144_sva_dfm_4_5 <= rva_out_reg_data_159_144_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_143_128_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_221_enex5 ) begin
      rva_out_reg_data_143_128_sva_dfm_4_5 <= rva_out_reg_data_143_128_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_222_enex5 ) begin
      rva_out_reg_data_127_112_sva_dfm_4_5 <= rva_out_reg_data_127_112_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_96_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_223_enex5 ) begin
      rva_out_reg_data_111_96_sva_dfm_4_5 <= rva_out_reg_data_111_96_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_80_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_224_enex5 ) begin
      rva_out_reg_data_95_80_sva_dfm_4_5 <= rva_out_reg_data_95_80_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_4_5 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_225_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_4_5 <= rva_out_reg_data_79_64_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_36_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_68_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_37_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_69_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_39_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_71_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1
          <= 16'b0000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[255:240]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_234_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[255:240]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_249_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[255:240]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_174_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_63_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[255:240]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_189_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_79_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[255:240]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_204_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_95_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[255:240]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_219_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[239:224]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_235_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[239:224]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_250_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[239:224]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_175_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[239:224]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_190_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_78_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[239:224]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_205_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_94_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[239:224]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_220_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[223:208]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_236_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[223:208]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_251_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[223:208]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_176_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_61_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[223:208]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_191_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_77_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[223:208]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_206_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_93_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[223:208]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_221_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[207:192]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_237_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[207:192]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_252_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[207:192]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_177_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_60_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[207:192]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_192_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_76_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[207:192]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_207_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_92_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[207:192]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_222_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_238_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_20_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_253_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_36_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_178_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_52_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_193_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_68_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_208_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_84_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[79:64]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_223_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[191:176]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_239_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[191:176]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_254_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[191:176]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_179_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_59_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[191:176]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_194_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_75_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[191:176]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_209_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_91_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[191:176]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_224_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_240_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_255_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_37_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_180_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_53_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_195_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_69_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_210_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_85_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[95:80]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_225_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[175:160]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_241_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[175:160]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[175:160]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_181_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_58_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[175:160]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_196_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_74_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[175:160]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_211_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_90_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[175:160]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_226_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_242_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_257_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_182_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_197_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_70_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_212_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_86_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[111:96]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_227_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_9_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[159:144]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_243_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[159:144]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[159:144]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_183_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_57_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[159:144]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_198_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_73_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[159:144]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_213_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_89_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[159:144]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_228_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_244_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_259_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_39_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_184_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_55_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_199_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_71_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_214_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_87_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[127:112]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_229_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_8_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[143:128]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_245_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[143:128]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_260_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[143:128]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_185_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_56_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[143:128]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_200_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_72_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[143:128]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_215_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_88_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[143:128]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_230_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6 <= 2'b00;
    end
    else if ( PECoreRun_wen & (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1
        | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1
        | and_dcpl_253) & and_dcpl_56 ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_3_7_6 <= weight_mem_write_arbxbar_xbar_for_empty_sva_2[7:6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1
          <= 16'b0000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_72_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[63:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_246_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[47:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_247_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1
          <= 16'b0000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_73_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_19_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, mux1h_2_nl, not_2436_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_18_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, mux1h_3_nl, not_2438_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, mux1h_4_nl, not_2440_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1
          <= 16'b0000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_74_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_51_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[63:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_201_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_50_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[47:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_202_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[31:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_203_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1
          <= 16'b0000000000000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1
          <= 16'b0000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_75_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_83_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[63:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_231_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[31:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_233_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1
        & while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_82_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[47:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_232_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_258 & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]))
        & nor_335_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[15:0]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_140_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1
          <= 16'b0000000000000000;
    end
    else if ( PECoreRun_wen & (~ mux_49_nl) & while_stage_0_6 ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_16_itm_1
          <= MUX_v_16_2_2(16'b0000000000000000, mux_348_nl, nand_67_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_1
          <= 1'b0;
    end
    else if ( weight_read_addrs_and_23_cse ) begin
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= weight_read_addrs_3_lpi_1_dfm_1[2:0];
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_31_itm_1
          <= ~((weight_read_addrs_3_lpi_1_dfm_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_data_sva_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rva_in_reg_data_and_tmp ) begin
      rva_in_reg_data_sva_1 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_284 & while_stage_0_7 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]))) & while_stage_0_4 )
        begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_9 <= 1'b0;
      rva_in_reg_rw_sva_st_9 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_9_cse ) begin
      rva_in_reg_rw_sva_st_1_9 <= rva_in_reg_rw_sva_st_1_8;
      rva_in_reg_rw_sva_st_9 <= rva_in_reg_rw_sva_st_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_1 <= 1'b0;
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( pe_manager_base_weight_and_5_cse ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_16_itm_1 <= pe_manager_base_weight_sva[0];
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_396_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_263_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_262_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_398_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_135_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_134_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_132_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_31_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_402_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= MUX_v_3_2_2((weight_read_addrs_1_lpi_1_dfm_1[2:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse
        & and_dcpl_274 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_15_itm_1
          <= ~((weight_read_addrs_1_lpi_1_dfm_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_159_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_359_itm_1
          & (pe_manager_base_weight_sva[1:0]==2'b11) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b110)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b101)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_1
          <= ~((pe_manager_base_weight_sva[2:0]!=3'b000));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_8_itm_1
          <= ~(pe_manager_base_weight_slc_pe_manager_base_weight_2_0_359_itm_1 |
          (pe_manager_base_weight_sva[1:0]!=2'b00));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_59_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_mx0w0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_52_itm_1 <= (pe_manager_base_weight_sva[2])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_153_itm_1 & (pe_manager_base_weight_sva[0])
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_48_itm_1 <= (pe_manager_base_weight_sva[1])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_141_itm_1 & (~
          (pe_manager_base_weight_sva[2])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_42_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_359_itm_1
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_141_itm_1 & (~
          (pe_manager_base_weight_sva[1])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1 <= (pe_manager_base_weight_sva[1])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_141_itm_1 & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1 <= (pe_manager_base_weight_sva[2])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_153_itm_1 & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_5_itm_1
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= (pe_manager_base_weight_sva[2])
          & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_4_itm_1
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1 <= (pe_manager_base_weight_sva[1:0]==2'b11)
          & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1 & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_1_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_8_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_153_itm_1
          & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_6_itm_1
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_163_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_nl,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_40_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1,
          PECore_UpdateFSM_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_mx0w0,
          PECore_RunFSM_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_50_nl & while_stage_0_5 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          input_read_req_valid_lpi_1_dfm_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_18_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_4 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_4 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_65_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_66_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_67_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_68_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_18_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_53_nl) & while_stage_0_5 ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= MUX_s_1_2_2((weight_read_addrs_4_14_2_lpi_1_dfm_1[0]),
          weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_9 <= 1'b0;
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_ftd <= 2'b00;
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_ftd_1 <= 2'b00;
      rva_out_reg_data_47_sva_dfm_4_4 <= 1'b0;
      rva_out_reg_data_63_sva_dfm_4_4 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( input_read_req_valid_and_2_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_9 <= input_read_req_valid_lpi_1_dfm_1_8;
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_ftd <= rva_out_reg_data_35_32_sva_dfm_4_3_rsp_0;
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_35_32_sva_dfm_4_3_rsp_1;
      rva_out_reg_data_47_sva_dfm_4_4 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      rva_out_reg_data_63_sva_dfm_4_4 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_11_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_7_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_226_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_7_1 <= rva_out_reg_data_23_17_sva_dfm_6_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_227_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= rva_out_reg_data_15_9_sva_dfm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_4 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_205_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_4 <= weight_port_read_out_data_0_0_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_228_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_4 <= rva_out_reg_data_39_36_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_229_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_4 <= rva_out_reg_data_46_40_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_4_4 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_230_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_4_4 <= rva_out_reg_data_62_48_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_255_240_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_231_enex5 ) begin
      rva_out_reg_data_255_240_sva_dfm_4_4 <= rva_out_reg_data_255_240_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_239_224_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_232_enex5 ) begin
      rva_out_reg_data_239_224_sva_dfm_4_4 <= rva_out_reg_data_239_224_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_223_208_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_233_enex5 ) begin
      rva_out_reg_data_223_208_sva_dfm_4_4 <= rva_out_reg_data_223_208_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_207_192_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_234_enex5 ) begin
      rva_out_reg_data_207_192_sva_dfm_4_4 <= rva_out_reg_data_207_192_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_191_176_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_235_enex5 ) begin
      rva_out_reg_data_191_176_sva_dfm_4_4 <= rva_out_reg_data_191_176_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_175_160_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_236_enex5 ) begin
      rva_out_reg_data_175_160_sva_dfm_4_4 <= rva_out_reg_data_175_160_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_159_144_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_237_enex5 ) begin
      rva_out_reg_data_159_144_sva_dfm_4_4 <= rva_out_reg_data_159_144_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_143_128_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_238_enex5 ) begin
      rva_out_reg_data_143_128_sva_dfm_4_4 <= rva_out_reg_data_143_128_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_239_enex5 ) begin
      rva_out_reg_data_127_112_sva_dfm_4_4 <= rva_out_reg_data_127_112_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_96_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_240_enex5 ) begin
      rva_out_reg_data_111_96_sva_dfm_4_4 <= rva_out_reg_data_111_96_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_80_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_241_enex5 ) begin
      rva_out_reg_data_95_80_sva_dfm_4_4 <= rva_out_reg_data_95_80_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_4_4 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_242_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_4_4 <= rva_out_reg_data_79_64_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= 8'b00000000;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_empty_and_3_enex5 ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= weight_mem_write_arbxbar_xbar_for_empty_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_380_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]))) & while_stage_0_4 )
        begin
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_380_itm_1 <= MUX_s_1_2_2((pe_manager_base_weight_sva_mx1_3_0[1]),
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_57 & (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse)
        ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_8_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_8 <= 1'b0;
      rva_in_reg_rw_sva_st_8 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_12_cse ) begin
      rva_in_reg_rw_sva_st_1_8 <= rva_in_reg_rw_sva_st_1_7;
      rva_in_reg_rw_sva_st_8 <= rva_in_reg_rw_sva_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_27_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_69_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_70_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_71_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_72_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_1_1_15 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_128_ssc ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
      weight_port_read_out_data_0_1_sva_dfm_1_1_15 <= MUX1HOT_s_1_9_2(weight_port_read_out_data_0_1_sva_mx0_15,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[31]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[15]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
          , weight_mem_run_3_for_5_and_158_ssc , weight_mem_run_3_for_5_and_159_ssc
          , weight_mem_run_3_for_5_and_160_ssc , weight_mem_run_3_for_5_and_161_ssc
          , weight_mem_run_3_for_5_and_162_cse , weight_mem_run_3_for_5_and_163_cse
          , weight_mem_run_3_for_5_and_164_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= MUX_v_256_256_2(input_mem_banks_bank_a_0_sva_dfm_2,
          input_mem_banks_bank_a_1_sva_dfm_2, input_mem_banks_bank_a_2_sva_dfm_2,
          input_mem_banks_bank_a_3_sva_dfm_2, input_mem_banks_bank_a_4_sva_dfm_2,
          input_mem_banks_bank_a_5_sva_dfm_2, input_mem_banks_bank_a_6_sva_dfm_2,
          input_mem_banks_bank_a_7_sva_dfm_2, input_mem_banks_bank_a_8_sva_dfm_2,
          input_mem_banks_bank_a_9_sva_dfm_2, input_mem_banks_bank_a_10_sva_dfm_2,
          input_mem_banks_bank_a_11_sva_dfm_2, input_mem_banks_bank_a_12_sva_dfm_2,
          input_mem_banks_bank_a_13_sva_dfm_2, input_mem_banks_bank_a_14_sva_dfm_2,
          input_mem_banks_bank_a_15_sva_dfm_2, input_mem_banks_bank_a_16_sva_dfm_2,
          input_mem_banks_bank_a_17_sva_dfm_2, input_mem_banks_bank_a_18_sva_dfm_2,
          input_mem_banks_bank_a_19_sva_dfm_2, input_mem_banks_bank_a_20_sva_dfm_2,
          input_mem_banks_bank_a_21_sva_dfm_2, input_mem_banks_bank_a_22_sva_dfm_2,
          input_mem_banks_bank_a_23_sva_dfm_2, input_mem_banks_bank_a_24_sva_dfm_2,
          input_mem_banks_bank_a_25_sva_dfm_2, input_mem_banks_bank_a_26_sva_dfm_2,
          input_mem_banks_bank_a_27_sva_dfm_2, input_mem_banks_bank_a_28_sva_dfm_2,
          input_mem_banks_bank_a_29_sva_dfm_2, input_mem_banks_bank_a_30_sva_dfm_2,
          input_mem_banks_bank_a_31_sva_dfm_2, input_mem_banks_bank_a_32_sva_dfm_2,
          input_mem_banks_bank_a_33_sva_dfm_2, input_mem_banks_bank_a_34_sva_dfm_2,
          input_mem_banks_bank_a_35_sva_dfm_2, input_mem_banks_bank_a_36_sva_dfm_2,
          input_mem_banks_bank_a_37_sva_dfm_2, input_mem_banks_bank_a_38_sva_dfm_2,
          input_mem_banks_bank_a_39_sva_dfm_2, input_mem_banks_bank_a_40_sva_dfm_2,
          input_mem_banks_bank_a_41_sva_dfm_2, input_mem_banks_bank_a_42_sva_dfm_2,
          input_mem_banks_bank_a_43_sva_dfm_2, input_mem_banks_bank_a_44_sva_dfm_2,
          input_mem_banks_bank_a_45_sva_dfm_2, input_mem_banks_bank_a_46_sva_dfm_2,
          input_mem_banks_bank_a_47_sva_dfm_2, input_mem_banks_bank_a_48_sva_dfm_2,
          input_mem_banks_bank_a_49_sva_dfm_2, input_mem_banks_bank_a_50_sva_dfm_2,
          input_mem_banks_bank_a_51_sva_dfm_2, input_mem_banks_bank_a_52_sva_dfm_2,
          input_mem_banks_bank_a_53_sva_dfm_2, input_mem_banks_bank_a_54_sva_dfm_2,
          input_mem_banks_bank_a_55_sva_dfm_2, input_mem_banks_bank_a_56_sva_dfm_2,
          input_mem_banks_bank_a_57_sva_dfm_2, input_mem_banks_bank_a_58_sva_dfm_2,
          input_mem_banks_bank_a_59_sva_dfm_2, input_mem_banks_bank_a_60_sva_dfm_2,
          input_mem_banks_bank_a_61_sva_dfm_2, input_mem_banks_bank_a_62_sva_dfm_2,
          input_mem_banks_bank_a_63_sva_dfm_2, input_mem_banks_bank_a_64_sva_dfm_2,
          input_mem_banks_bank_a_65_sva_dfm_2, input_mem_banks_bank_a_66_sva_dfm_2,
          input_mem_banks_bank_a_67_sva_dfm_2, input_mem_banks_bank_a_68_sva_dfm_2,
          input_mem_banks_bank_a_69_sva_dfm_2, input_mem_banks_bank_a_70_sva_dfm_2,
          input_mem_banks_bank_a_71_sva_dfm_2, input_mem_banks_bank_a_72_sva_dfm_2,
          input_mem_banks_bank_a_73_sva_dfm_2, input_mem_banks_bank_a_74_sva_dfm_2,
          input_mem_banks_bank_a_75_sva_dfm_2, input_mem_banks_bank_a_76_sva_dfm_2,
          input_mem_banks_bank_a_77_sva_dfm_2, input_mem_banks_bank_a_78_sva_dfm_2,
          input_mem_banks_bank_a_79_sva_dfm_2, input_mem_banks_bank_a_80_sva_dfm_2,
          input_mem_banks_bank_a_81_sva_dfm_2, input_mem_banks_bank_a_82_sva_dfm_2,
          input_mem_banks_bank_a_83_sva_dfm_2, input_mem_banks_bank_a_84_sva_dfm_2,
          input_mem_banks_bank_a_85_sva_dfm_2, input_mem_banks_bank_a_86_sva_dfm_2,
          input_mem_banks_bank_a_87_sva_dfm_2, input_mem_banks_bank_a_88_sva_dfm_2,
          input_mem_banks_bank_a_89_sva_dfm_2, input_mem_banks_bank_a_90_sva_dfm_2,
          input_mem_banks_bank_a_91_sva_dfm_2, input_mem_banks_bank_a_92_sva_dfm_2,
          input_mem_banks_bank_a_93_sva_dfm_2, input_mem_banks_bank_a_94_sva_dfm_2,
          input_mem_banks_bank_a_95_sva_dfm_2, input_mem_banks_bank_a_96_sva_dfm_2,
          input_mem_banks_bank_a_97_sva_dfm_2, input_mem_banks_bank_a_98_sva_dfm_2,
          input_mem_banks_bank_a_99_sva_dfm_2, input_mem_banks_bank_a_100_sva_dfm_2,
          input_mem_banks_bank_a_101_sva_dfm_2, input_mem_banks_bank_a_102_sva_dfm_2,
          input_mem_banks_bank_a_103_sva_dfm_2, input_mem_banks_bank_a_104_sva_dfm_2,
          input_mem_banks_bank_a_105_sva_dfm_2, input_mem_banks_bank_a_106_sva_dfm_2,
          input_mem_banks_bank_a_107_sva_dfm_2, input_mem_banks_bank_a_108_sva_dfm_2,
          input_mem_banks_bank_a_109_sva_dfm_2, input_mem_banks_bank_a_110_sva_dfm_2,
          input_mem_banks_bank_a_111_sva_dfm_2, input_mem_banks_bank_a_112_sva_dfm_2,
          input_mem_banks_bank_a_113_sva_dfm_2, input_mem_banks_bank_a_114_sva_dfm_2,
          input_mem_banks_bank_a_115_sva_dfm_2, input_mem_banks_bank_a_116_sva_dfm_2,
          input_mem_banks_bank_a_117_sva_dfm_2, input_mem_banks_bank_a_118_sva_dfm_2,
          input_mem_banks_bank_a_119_sva_dfm_2, input_mem_banks_bank_a_120_sva_dfm_2,
          input_mem_banks_bank_a_121_sva_dfm_2, input_mem_banks_bank_a_122_sva_dfm_2,
          input_mem_banks_bank_a_123_sva_dfm_2, input_mem_banks_bank_a_124_sva_dfm_2,
          input_mem_banks_bank_a_125_sva_dfm_2, input_mem_banks_bank_a_126_sva_dfm_2,
          input_mem_banks_bank_a_127_sva_dfm_2, input_mem_banks_bank_a_128_sva_dfm_2,
          input_mem_banks_bank_a_129_sva_dfm_2, input_mem_banks_bank_a_130_sva_dfm_2,
          input_mem_banks_bank_a_131_sva_dfm_2, input_mem_banks_bank_a_132_sva_dfm_2,
          input_mem_banks_bank_a_133_sva_dfm_2, input_mem_banks_bank_a_134_sva_dfm_2,
          input_mem_banks_bank_a_135_sva_dfm_2, input_mem_banks_bank_a_136_sva_dfm_2,
          input_mem_banks_bank_a_137_sva_dfm_2, input_mem_banks_bank_a_138_sva_dfm_2,
          input_mem_banks_bank_a_139_sva_dfm_2, input_mem_banks_bank_a_140_sva_dfm_2,
          input_mem_banks_bank_a_141_sva_dfm_2, input_mem_banks_bank_a_142_sva_dfm_2,
          input_mem_banks_bank_a_143_sva_dfm_2, input_mem_banks_bank_a_144_sva_dfm_2,
          input_mem_banks_bank_a_145_sva_dfm_2, input_mem_banks_bank_a_146_sva_dfm_2,
          input_mem_banks_bank_a_147_sva_dfm_2, input_mem_banks_bank_a_148_sva_dfm_2,
          input_mem_banks_bank_a_149_sva_dfm_2, input_mem_banks_bank_a_150_sva_dfm_2,
          input_mem_banks_bank_a_151_sva_dfm_2, input_mem_banks_bank_a_152_sva_dfm_2,
          input_mem_banks_bank_a_153_sva_dfm_2, input_mem_banks_bank_a_154_sva_dfm_2,
          input_mem_banks_bank_a_155_sva_dfm_2, input_mem_banks_bank_a_156_sva_dfm_2,
          input_mem_banks_bank_a_157_sva_dfm_2, input_mem_banks_bank_a_158_sva_dfm_2,
          input_mem_banks_bank_a_159_sva_dfm_2, input_mem_banks_bank_a_160_sva_dfm_2,
          input_mem_banks_bank_a_161_sva_dfm_2, input_mem_banks_bank_a_162_sva_dfm_2,
          input_mem_banks_bank_a_163_sva_dfm_2, input_mem_banks_bank_a_164_sva_dfm_2,
          input_mem_banks_bank_a_165_sva_dfm_2, input_mem_banks_bank_a_166_sva_dfm_2,
          input_mem_banks_bank_a_167_sva_dfm_2, input_mem_banks_bank_a_168_sva_dfm_2,
          input_mem_banks_bank_a_169_sva_dfm_2, input_mem_banks_bank_a_170_sva_dfm_2,
          input_mem_banks_bank_a_171_sva_dfm_2, input_mem_banks_bank_a_172_sva_dfm_2,
          input_mem_banks_bank_a_173_sva_dfm_2, input_mem_banks_bank_a_174_sva_dfm_2,
          input_mem_banks_bank_a_175_sva_dfm_2, input_mem_banks_bank_a_176_sva_dfm_2,
          input_mem_banks_bank_a_177_sva_dfm_2, input_mem_banks_bank_a_178_sva_dfm_2,
          input_mem_banks_bank_a_179_sva_dfm_2, input_mem_banks_bank_a_180_sva_dfm_2,
          input_mem_banks_bank_a_181_sva_dfm_2, input_mem_banks_bank_a_182_sva_dfm_2,
          input_mem_banks_bank_a_183_sva_dfm_2, input_mem_banks_bank_a_184_sva_dfm_2,
          input_mem_banks_bank_a_185_sva_dfm_2, input_mem_banks_bank_a_186_sva_dfm_2,
          input_mem_banks_bank_a_187_sva_dfm_2, input_mem_banks_bank_a_188_sva_dfm_2,
          input_mem_banks_bank_a_189_sva_dfm_2, input_mem_banks_bank_a_190_sva_dfm_2,
          input_mem_banks_bank_a_191_sva_dfm_2, input_mem_banks_bank_a_192_sva_dfm_2,
          input_mem_banks_bank_a_193_sva_dfm_2, input_mem_banks_bank_a_194_sva_dfm_2,
          input_mem_banks_bank_a_195_sva_dfm_2, input_mem_banks_bank_a_196_sva_dfm_2,
          input_mem_banks_bank_a_197_sva_dfm_2, input_mem_banks_bank_a_198_sva_dfm_2,
          input_mem_banks_bank_a_199_sva_dfm_2, input_mem_banks_bank_a_200_sva_dfm_2,
          input_mem_banks_bank_a_201_sva_dfm_2, input_mem_banks_bank_a_202_sva_dfm_2,
          input_mem_banks_bank_a_203_sva_dfm_2, input_mem_banks_bank_a_204_sva_dfm_2,
          input_mem_banks_bank_a_205_sva_dfm_2, input_mem_banks_bank_a_206_sva_dfm_2,
          input_mem_banks_bank_a_207_sva_dfm_2, input_mem_banks_bank_a_208_sva_dfm_2,
          input_mem_banks_bank_a_209_sva_dfm_2, input_mem_banks_bank_a_210_sva_dfm_2,
          input_mem_banks_bank_a_211_sva_dfm_2, input_mem_banks_bank_a_212_sva_dfm_2,
          input_mem_banks_bank_a_213_sva_dfm_2, input_mem_banks_bank_a_214_sva_dfm_2,
          input_mem_banks_bank_a_215_sva_dfm_2, input_mem_banks_bank_a_216_sva_dfm_2,
          input_mem_banks_bank_a_217_sva_dfm_2, input_mem_banks_bank_a_218_sva_dfm_2,
          input_mem_banks_bank_a_219_sva_dfm_2, input_mem_banks_bank_a_220_sva_dfm_2,
          input_mem_banks_bank_a_221_sva_dfm_2, input_mem_banks_bank_a_222_sva_dfm_2,
          input_mem_banks_bank_a_223_sva_dfm_2, input_mem_banks_bank_a_224_sva_dfm_2,
          input_mem_banks_bank_a_225_sva_dfm_2, input_mem_banks_bank_a_226_sva_dfm_2,
          input_mem_banks_bank_a_227_sva_dfm_2, input_mem_banks_bank_a_228_sva_dfm_2,
          input_mem_banks_bank_a_229_sva_dfm_2, input_mem_banks_bank_a_230_sva_dfm_2,
          input_mem_banks_bank_a_231_sva_dfm_2, input_mem_banks_bank_a_232_sva_dfm_2,
          input_mem_banks_bank_a_233_sva_dfm_2, input_mem_banks_bank_a_234_sva_dfm_2,
          input_mem_banks_bank_a_235_sva_dfm_2, input_mem_banks_bank_a_236_sva_dfm_2,
          input_mem_banks_bank_a_237_sva_dfm_2, input_mem_banks_bank_a_238_sva_dfm_2,
          input_mem_banks_bank_a_239_sva_dfm_2, input_mem_banks_bank_a_240_sva_dfm_2,
          input_mem_banks_bank_a_241_sva_dfm_2, input_mem_banks_bank_a_242_sva_dfm_2,
          input_mem_banks_bank_a_243_sva_dfm_2, input_mem_banks_bank_a_244_sva_dfm_2,
          input_mem_banks_bank_a_245_sva_dfm_2, input_mem_banks_bank_a_246_sva_dfm_2,
          input_mem_banks_bank_a_247_sva_dfm_2, input_mem_banks_bank_a_248_sva_dfm_2,
          input_mem_banks_bank_a_249_sva_dfm_2, input_mem_banks_bank_a_250_sva_dfm_2,
          input_mem_banks_bank_a_251_sva_dfm_2, input_mem_banks_bank_a_252_sva_dfm_2,
          input_mem_banks_bank_a_253_sva_dfm_2, input_mem_banks_bank_a_254_sva_dfm_2,
          input_mem_banks_bank_a_255_sva_dfm_2, input_mem_banks_read_1_for_mux_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= 1'b0;
      rva_out_reg_data_35_32_sva_dfm_4_3_rsp_0 <= 2'b00;
      rva_out_reg_data_35_32_sva_dfm_4_3_rsp_1 <= 2'b00;
    end
    else if ( input_read_req_valid_and_3_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= input_read_req_valid_lpi_1_dfm_1_7;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
      rva_out_reg_data_35_32_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_35_32_sva_dfm_4_2_3_2;
      rva_out_reg_data_35_32_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_35_32_sva_dfm_4_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_15_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_6_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_243_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_6_1 <= rva_out_reg_data_23_17_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_244_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= rva_out_reg_data_15_9_sva_dfm_7_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_3 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_206_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_3 <= weight_port_read_out_data_0_0_sva_dfm_2_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_168_cse ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd <= weight_port_read_out_data_0_1_sva_dfm_2_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_207_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1 <= weight_port_read_out_data_0_1_sva_dfm_2_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_245_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_3 <= rva_out_reg_data_39_36_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_246_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3 <= rva_out_reg_data_46_40_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_4_3 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_247_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_4_3 <= rva_out_reg_data_62_48_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_255_240_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_248_enex5 ) begin
      rva_out_reg_data_255_240_sva_dfm_4_3 <= rva_out_reg_data_255_240_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_239_224_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_249_enex5 ) begin
      rva_out_reg_data_239_224_sva_dfm_4_3 <= rva_out_reg_data_239_224_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_223_208_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_250_enex5 ) begin
      rva_out_reg_data_223_208_sva_dfm_4_3 <= rva_out_reg_data_223_208_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_207_192_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_251_enex5 ) begin
      rva_out_reg_data_207_192_sva_dfm_4_3 <= rva_out_reg_data_207_192_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_191_176_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_252_enex5 ) begin
      rva_out_reg_data_191_176_sva_dfm_4_3 <= rva_out_reg_data_191_176_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_175_160_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_253_enex5 ) begin
      rva_out_reg_data_175_160_sva_dfm_4_3 <= rva_out_reg_data_175_160_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_159_144_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_254_enex5 ) begin
      rva_out_reg_data_159_144_sva_dfm_4_3 <= rva_out_reg_data_159_144_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_143_128_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_255_enex5 ) begin
      rva_out_reg_data_143_128_sva_dfm_4_3 <= rva_out_reg_data_143_128_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_256_enex5 ) begin
      rva_out_reg_data_127_112_sva_dfm_4_3 <= rva_out_reg_data_127_112_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_96_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_257_enex5 ) begin
      rva_out_reg_data_111_96_sva_dfm_4_3 <= rva_out_reg_data_111_96_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_80_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_258_enex5 ) begin
      rva_out_reg_data_95_80_sva_dfm_4_3 <= rva_out_reg_data_95_80_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_4_3 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_259_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_4_3 <= rva_out_reg_data_79_64_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_234_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_182)
        ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_234_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_238_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_189)
        ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_238_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_242_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_193)
        ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_242_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_246_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_197)
        ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_246_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_250_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_201)
        ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_250_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_254_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_203)
        ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_254_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_258_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_205)
        ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_258_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_262_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_207)
        ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_262_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_266_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_211)
        ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_266_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_270_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_213)
        ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_270_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_274_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_215)
        ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_274_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_278_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_217)
        ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_278_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_282_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_221)
        ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_282_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_286_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_223)
        ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_286_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_290_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_225)
        ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_290_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_294_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_227)
        ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_294_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_298_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_230)
        ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_298_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_302_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_232)
        ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_302_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_306_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_234)
        ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_306_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_310_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_236)
        ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_310_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_314_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_239)
        ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_314_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_318_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_241)
        ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_318_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_322_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_243)
        ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_322_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_326_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_245)
        ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_326_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_330_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_248)
        ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_330_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_334_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_250)
        ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_334_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_338_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_252)
        ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_338_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_342_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_254)
        ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_342_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_346_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_257)
        ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_346_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_350_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_259)
        ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_350_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_354_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_261)
        ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_354_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_358_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_263)
        ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_358_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_362_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_267)
        ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_362_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_366_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_270)
        ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_366_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_370_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_273)
        ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_370_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_374_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_276)
        ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_374_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_378_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_278)
        ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_378_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_382_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_280)
        ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_382_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_386_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_282)
        ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_386_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_390_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_284)
        ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_390_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_394_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_286)
        ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_394_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_398_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_288)
        ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_398_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_402_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_290)
        ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_402_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_406_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_292)
        ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_406_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_410_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_294)
        ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_410_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_414_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_296)
        ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_414_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_418_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_298)
        ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_418_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_422_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_300)
        ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_422_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_426_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_302)
        ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_426_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_430_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_304)
        ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_430_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_434_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_306)
        ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_434_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_438_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_308)
        ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_438_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_442_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_310)
        ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_442_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_446_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_312)
        ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_446_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_450_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_314)
        ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_450_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_454_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_316)
        ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_454_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_458_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_318)
        ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_458_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_462_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_320)
        ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_462_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_466_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_322)
        ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_466_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_470_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_324)
        ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_470_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_474_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_326)
        ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_474_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_478_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_328)
        ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_478_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_482_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_330)
        ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_482_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_486_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_332)
        ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_486_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_490_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_182)
        ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_490_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_494_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_189)
        ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_494_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_498_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_193)
        ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_498_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_502_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_197)
        ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_502_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_506_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_201)
        ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_506_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_510_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_203)
        ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_510_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_514_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_205)
        ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_514_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_518_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_207)
        ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_518_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_522_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_211)
        ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_522_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_526_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_213)
        ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_526_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_530_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_215)
        ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_530_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_534_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_217)
        ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_534_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_538_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_221)
        ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_538_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_542_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_223)
        ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_542_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_546_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_225)
        ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_546_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_550_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_227)
        ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_550_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_554_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_230)
        ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_554_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_558_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_232)
        ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_558_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_562_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_234)
        ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_562_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_566_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_236)
        ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_566_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_570_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_239)
        ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_570_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_574_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_241)
        ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_574_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_578_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_243)
        ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_578_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_582_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_245)
        ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_582_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_586_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_248)
        ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_586_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_590_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_250)
        ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_590_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_594_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_252)
        ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_594_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_598_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_254)
        ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_598_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_602_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_257)
        ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_602_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_606_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_259)
        ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_606_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_610_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_261)
        ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_610_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_614_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_263)
        ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_614_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_618_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_267)
        ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_618_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_622_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_270)
        ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_622_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_626_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_273)
        ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_626_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_630_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_276)
        ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_630_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_634_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_278)
        ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_634_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_638_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_280)
        ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_638_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_642_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_282)
        ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_642_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_646_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_284)
        ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_646_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_650_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_286)
        ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_650_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_654_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_288)
        ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_654_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_658_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_290)
        ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_658_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_662_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_292)
        ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_662_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_666_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_294)
        ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_666_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_670_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_296)
        ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_670_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_674_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_298)
        ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_674_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_678_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_300)
        ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_678_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_682_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_302)
        ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_682_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_686_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_304)
        ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_686_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_690_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_306)
        ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_690_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_694_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_308)
        ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_694_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_698_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_310)
        ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_698_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_702_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_312)
        ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_702_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_706_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_314)
        ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_706_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_710_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_316)
        ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_710_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_714_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_318)
        ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_714_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_718_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_320)
        ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_718_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_722_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_322)
        ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_722_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_726_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_324)
        ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_726_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_730_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_326)
        ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_730_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_734_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_328)
        ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_734_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_738_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_330)
        ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_738_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
        & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_742_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_332)
        ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_742_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_746_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_403)
        ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_746_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_750_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_406)
        ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_750_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_754_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_409)
        ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_754_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_758_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_412)
        ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_758_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_762_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_414)
        ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_762_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_766_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_416)
        ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_766_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_770_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_418)
        ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_770_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_774_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_420)
        ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_774_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_778_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_422)
        ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_778_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_782_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_424)
        ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_782_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_786_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_426)
        ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_786_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_790_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_428)
        ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_790_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_794_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_430)
        ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_794_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_798_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_432)
        ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_798_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_802_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_434)
        ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_802_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_806_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_436)
        ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_806_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_810_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_438)
        ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_810_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_814_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_440)
        ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_814_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_818_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_442)
        ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_818_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_822_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_444)
        ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_822_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_826_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_446)
        ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_826_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_830_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_448)
        ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_830_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_834_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_450)
        ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_834_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_838_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_452)
        ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_838_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_842_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_454)
        ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_842_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_846_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_456)
        ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_846_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_850_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_458)
        ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_850_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_854_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_460)
        ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_854_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_858_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_462)
        ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_858_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_862_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_464)
        ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_862_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_866_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_466)
        ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_866_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_870_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_468)
        ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_870_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_874_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_472)
        ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_874_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_878_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_475)
        ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_878_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_882_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_478)
        ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_882_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_886_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_481)
        ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_886_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_890_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_483)
        ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_890_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_894_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_485)
        ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_894_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_898_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_487)
        ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_898_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_902_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_489)
        ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_902_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_906_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_491)
        ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_906_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_910_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_493)
        ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_910_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_914_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_495)
        ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_914_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_918_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_497)
        ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_918_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_922_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_499)
        ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_922_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_926_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_501)
        ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_926_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_930_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_503)
        ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_930_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_934_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_505)
        ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_934_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_938_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_507)
        ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_938_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_942_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_509)
        ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_942_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_946_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_511)
        ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_946_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_950_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_513)
        ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_950_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_954_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_515)
        ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_954_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_958_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_517)
        ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_958_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_962_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_519)
        ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_962_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_966_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_521)
        ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_966_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_970_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_523)
        ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_970_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_974_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_525)
        ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_974_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_978_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_527)
        ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_978_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_982_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_529)
        ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_982_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_986_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_531)
        ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_986_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_990_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_533)
        ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_990_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_994_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_535)
        ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_994_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_998_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_185 | or_dcpl_537)
        ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_998_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1002_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_403)
        ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1002_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1006_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_406)
        ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1006_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1010_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_409)
        ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1010_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1014_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_412)
        ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1014_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1018_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_414)
        ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1018_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1022_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_416)
        ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1022_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1026_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_418)
        ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1026_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1030_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_420)
        ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1030_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1034_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_422)
        ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1034_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1038_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_424)
        ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1038_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1042_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_426)
        ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1042_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1046_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_428)
        ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1046_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1050_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_430)
        ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1050_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1054_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_432)
        ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1054_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1058_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_434)
        ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1058_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1062_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_436)
        ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1062_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1066_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_438)
        ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1066_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1070_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_440)
        ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1070_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1074_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_442)
        ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1074_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1078_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_444)
        ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1078_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1082_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_446)
        ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1082_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1086_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_448)
        ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1086_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1090_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_450)
        ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1090_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1094_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_452)
        ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1094_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1098_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_454)
        ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1098_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1102_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_456)
        ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1102_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1106_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_458)
        ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1106_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1110_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_460)
        ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1110_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1114_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_462)
        ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1114_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1118_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_464)
        ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1118_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1122_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_466)
        ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1122_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1126_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_468)
        ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1126_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1130_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_472)
        ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1130_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1134_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_475)
        ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1134_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1138_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_478)
        ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1138_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1142_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_481)
        ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1142_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1146_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_483)
        ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1146_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1150_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_485)
        ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1150_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1154_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_487)
        ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1154_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1158_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_489)
        ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1158_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1162_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_491)
        ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1162_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1166_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_493)
        ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1166_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1170_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_495)
        ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1170_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1174_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_497)
        ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1174_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1178_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_499)
        ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1178_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1182_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_501)
        ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1182_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1186_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_503)
        ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1186_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1190_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_505)
        ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1190_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1194_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_507)
        ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1194_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1198_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_509)
        ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1198_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1202_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_511)
        ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1202_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1206_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_513)
        ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1206_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1210_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_515)
        ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1210_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1214_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_517)
        ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1214_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1218_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_519)
        ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1218_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1222_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_521)
        ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1222_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1226_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_523)
        ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1226_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1230_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_525)
        ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1230_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1234_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_527)
        ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1234_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1238_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_529)
        ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1238_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1242_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_531)
        ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1242_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1246_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_533)
        ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1246_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1250_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_535)
        ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1250_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & ((input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
        & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        | while_and_1254_rgt) & while_stage_0_3 & fsm_output & (or_dcpl_336 | or_dcpl_537)
        ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= MUX_v_256_2_2(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
          rva_in_reg_data_sva_1, while_and_1254_rgt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_7 <= 1'b0;
      rva_in_reg_rw_sva_st_7 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_15_cse ) begin
      rva_in_reg_rw_sva_st_1_7 <= rva_in_reg_rw_sva_st_1_6;
      rva_in_reg_rw_sva_st_7 <= rva_in_reg_rw_sva_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_36_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_73_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_74_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_75_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_76_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= 1'b0;
      rva_out_reg_data_35_32_sva_dfm_4_2_3_2 <= 2'b00;
      rva_out_reg_data_35_32_sva_dfm_4_2_1_0 <= 2'b00;
    end
    else if ( input_read_req_valid_and_4_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= input_read_req_valid_lpi_1_dfm_1_6;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
      rva_out_reg_data_35_32_sva_dfm_4_2_3_2 <= rva_out_reg_data_35_32_sva_dfm_4_1_3_2;
      rva_out_reg_data_35_32_sva_dfm_4_2_1_0 <= rva_out_reg_data_35_32_sva_dfm_4_1_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_19_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_ftd <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_260_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_ftd <= rva_out_reg_data_30_25_sva_dfm_4_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_ftd_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_108_ssc ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_ftd_1 <= rva_out_reg_data_30_25_sva_dfm_4_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_261_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= rva_out_reg_data_23_17_sva_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_7_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_262_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_7_1 <= rva_out_reg_data_15_9_sva_dfm_6_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_1 <= 16'b0000000000000000;
    end
    else if ( weight_port_read_out_data_and_208_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_1 <= weight_port_read_out_data_0_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_263_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_4_2 <= rva_out_reg_data_39_36_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_264_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2 <= rva_out_reg_data_46_40_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_4_2 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_265_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_4_2 <= rva_out_reg_data_62_48_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_255_240_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_266_enex5 ) begin
      rva_out_reg_data_255_240_sva_dfm_4_2 <= rva_out_reg_data_255_240_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_239_224_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_267_enex5 ) begin
      rva_out_reg_data_239_224_sva_dfm_4_2 <= rva_out_reg_data_239_224_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_223_208_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_268_enex5 ) begin
      rva_out_reg_data_223_208_sva_dfm_4_2 <= rva_out_reg_data_223_208_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_207_192_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_269_enex5 ) begin
      rva_out_reg_data_207_192_sva_dfm_4_2 <= rva_out_reg_data_207_192_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_191_176_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_270_enex5 ) begin
      rva_out_reg_data_191_176_sva_dfm_4_2 <= rva_out_reg_data_191_176_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_175_160_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_271_enex5 ) begin
      rva_out_reg_data_175_160_sva_dfm_4_2 <= rva_out_reg_data_175_160_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_159_144_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_272_enex5 ) begin
      rva_out_reg_data_159_144_sva_dfm_4_2 <= rva_out_reg_data_159_144_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_143_128_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_273_enex5 ) begin
      rva_out_reg_data_143_128_sva_dfm_4_2 <= rva_out_reg_data_143_128_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_127_112_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_274_enex5 ) begin
      rva_out_reg_data_127_112_sva_dfm_4_2 <= rva_out_reg_data_127_112_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_111_96_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_275_enex5 ) begin
      rva_out_reg_data_111_96_sva_dfm_4_2 <= rva_out_reg_data_111_96_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_95_80_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_276_enex5 ) begin
      rva_out_reg_data_95_80_sva_dfm_4_2 <= rva_out_reg_data_95_80_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_4_2 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_277_enex5 ) begin
      rva_out_reg_data_79_64_sva_dfm_4_2 <= rva_out_reg_data_79_64_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_base_input_and_tmp ) begin
      pe_manager_base_input_sva <= MUX_v_15_2_2(pe_manager_base_input_sva_dfm_3_1,
          PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl,
          and_dcpl_180);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( (~((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01) & rva_in_PopNB_mioi_return_rsc_z_mxwt
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5:3]!=3'b000)))
        & nor_534_cse & nor_518_cse & nor_520_cse & nor_521_cse & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
        & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt))
        & while_stage_0_3)) & rva_in_reg_rw_and_4_cse ) begin
      pe_manager_base_input_sva_dfm_3_1 <= MUX_v_15_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[62:48]),
          pe_manager_base_input_sva_mx1, or_834_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_54_nl) & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_6 <= 1'b0;
      rva_in_reg_rw_sva_st_6 <= 1'b0;
      PECore_PushAxiRsp_mux_26_itm_1 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_1_15 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_131_cse ) begin
      rva_in_reg_rw_sva_st_1_6 <= rva_in_reg_rw_sva_st_1_5;
      rva_in_reg_rw_sva_st_6 <= rva_in_reg_rw_sva_st_5;
      PECore_PushAxiRsp_mux_26_itm_1 <= MUX_s_1_2_2(weight_port_read_out_data_mux_67_nl,
          rva_out_reg_data_63_sva_dfm_7, rva_in_reg_rw_sva_5);
      weight_port_read_out_data_0_1_sva_dfm_1_15 <= mux1h_1_nl & (~ or_dcpl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_45_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_4[0];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_4[8];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[16];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[31];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_77_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_78_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:9];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_79_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:17];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_80_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[30:25];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( input_read_req_valid_and_5_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_324_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_23_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_278_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_4 <= rva_out_reg_data_23_17_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_6_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_279_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_6_1 <= rva_out_reg_data_15_9_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_4_1 <= 7'b0000000;
      rva_out_reg_data_62_48_sva_dfm_4_1 <= 15'b000000000000000;
    end
    else if ( and_1344_cse ) begin
      rva_out_reg_data_39_36_sva_dfm_4_1 <= MUX1HOT_v_4_4_2(rva_out_reg_data_39_36_sva_dfm_1_5,
          rva_out_reg_data_39_36_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:36]),
          (weight_port_read_out_data_0_2_sva_dfm_2[7:4]), {PECore_PushAxiRsp_if_asn_93
          , PECore_PushAxiRsp_if_asn_95 , PECore_PushAxiRsp_if_asn_91 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_46_40_sva_dfm_4_1 <= MUX1HOT_v_7_4_2(rva_out_reg_data_46_40_sva_dfm_1_5,
          rva_out_reg_data_46_40_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[46:40]),
          (weight_port_read_out_data_0_2_sva_dfm_2[14:8]), {PECore_PushAxiRsp_if_asn_93
          , PECore_PushAxiRsp_if_asn_95 , PECore_PushAxiRsp_if_asn_91 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_62_48_sva_dfm_4_1 <= MUX1HOT_v_15_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0,
          rva_out_reg_data_62_48_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[62:48]),
          (weight_port_read_out_data_0_3_sva_dfm_2[14:0]), {PECore_PushAxiRsp_if_asn_93
          , PECore_PushAxiRsp_if_asn_95 , PECore_PushAxiRsp_if_asn_91 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_255_240_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_239_224_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_223_208_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_207_192_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_191_176_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_175_160_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_159_144_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_143_128_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_127_112_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_111_96_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_95_80_sva_dfm_4_1 <= 16'b0000000000000000;
      rva_out_reg_data_79_64_sva_dfm_4_1 <= 16'b0000000000000000;
    end
    else if ( rva_out_reg_data_and_134_cse ) begin
      rva_out_reg_data_255_240_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_255_240_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_13_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_port_read_out_data_6_12_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
      rva_out_reg_data_239_224_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_239_224_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_12_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_port_read_out_data_6_11_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
      rva_out_reg_data_223_208_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_223_208_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_11_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_port_read_out_data_6_10_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
      rva_out_reg_data_207_192_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_207_192_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_10_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_port_read_out_data_6_9_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
      rva_out_reg_data_191_176_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_191_176_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_9_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000,
          weight_port_read_out_data_6_8_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
      rva_out_reg_data_175_160_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_175_160_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000,
          weight_port_read_out_data_6_7_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
      rva_out_reg_data_159_144_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_159_144_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000,
          weight_port_read_out_data_6_6_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
      rva_out_reg_data_143_128_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_143_128_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000,
          weight_port_read_out_data_6_5_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
      rva_out_reg_data_127_112_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_127_112_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0_000000,
          weight_port_read_out_data_6_4_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
      rva_out_reg_data_111_96_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_111_96_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000006,
          weight_port_read_out_data_0_10_sva_dfm_2, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1256_cse , while_while_nor_259_cse});
      rva_out_reg_data_95_80_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_95_80_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000007,
          weight_port_read_out_data_0_11_sva_dfm_2, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1256_cse , while_while_nor_259_cse});
      rva_out_reg_data_79_64_sva_dfm_4_1 <= MUX1HOT_v_16_3_2(rva_out_reg_data_79_64_sva_dfm_4_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_14_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_15_0000000,
          weight_port_read_out_data_6_13_sva_dfm_1, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , and_dcpl_674 , and_dcpl_675});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_63_sva_dfm_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ nand_72_cse) ) begin
      rva_out_reg_data_63_sva_dfm_6 <= PECore_PushAxiRsp_mux_26_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_6 <= 15'b000000000000000;
      rva_out_reg_data_46_40_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_39_36_sva_dfm_6 <= 4'b0000;
    end
    else if ( and_1357_cse ) begin
      rva_out_reg_data_62_48_sva_dfm_6 <= rva_out_reg_data_62_48_sva_dfm_6_mx1;
      rva_out_reg_data_46_40_sva_dfm_6 <= rva_out_reg_data_46_40_sva_dfm_6_mx1;
      rva_out_reg_data_39_36_sva_dfm_6 <= rva_out_reg_data_39_36_sva_dfm_6_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(rva_in_reg_rw_sva_5 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        | (~ while_stage_0_7))) ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          (weight_port_read_out_data_0_2_sva_dfm_2[15]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_54_tmp ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= MUX1HOT_v_256_3_2(input_mem_banks_read_read_data_lpi_1_dfm_1_3,
          weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d, weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1,
          {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          , and_688_nl , nor_463_nl});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_280_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_5 <= rva_out_reg_data_46_40_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_5 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_281_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_5 <= rva_out_reg_data_39_36_sva_dfm_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_79_64_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_95_80_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_111_96_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_127_112_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_143_128_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_159_144_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_175_160_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_191_176_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_207_192_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_223_208_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_239_224_sva_dfm_6 <= 16'b0000000000000000;
      rva_out_reg_data_255_240_sva_dfm_6 <= 16'b0000000000000000;
    end
    else if ( and_1372_cse ) begin
      rva_out_reg_data_79_64_sva_dfm_6 <= rva_out_reg_data_79_64_sva_dfm_4_mx0w0;
      rva_out_reg_data_95_80_sva_dfm_6 <= rva_out_reg_data_95_80_sva_dfm_4_mx0w0;
      rva_out_reg_data_111_96_sva_dfm_6 <= rva_out_reg_data_111_96_sva_dfm_4_mx0w0;
      rva_out_reg_data_127_112_sva_dfm_6 <= rva_out_reg_data_127_112_sva_dfm_4_mx0w0;
      rva_out_reg_data_143_128_sva_dfm_6 <= rva_out_reg_data_143_128_sva_dfm_4_mx0w0;
      rva_out_reg_data_159_144_sva_dfm_6 <= rva_out_reg_data_159_144_sva_dfm_4_mx0w0;
      rva_out_reg_data_175_160_sva_dfm_6 <= rva_out_reg_data_175_160_sva_dfm_4_mx0w0;
      rva_out_reg_data_191_176_sva_dfm_6 <= rva_out_reg_data_191_176_sva_dfm_4_mx0w0;
      rva_out_reg_data_207_192_sva_dfm_6 <= rva_out_reg_data_207_192_sva_dfm_4_mx0w0;
      rva_out_reg_data_223_208_sva_dfm_6 <= rva_out_reg_data_223_208_sva_dfm_4_mx0w0;
      rva_out_reg_data_239_224_sva_dfm_6 <= rva_out_reg_data_239_224_sva_dfm_4_mx0w0;
      rva_out_reg_data_255_240_sva_dfm_6 <= rva_out_reg_data_255_240_sva_dfm_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_24_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_27_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_278_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_271_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_264_itm_1_1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_282_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_3 <= rva_out_reg_data_23_17_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_283_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_5 <= rva_out_reg_data_15_9_sva_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_28_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= 1'b0;
      rva_out_reg_data_35_32_sva_dfm_1_4_3_2 <= 2'b00;
      rva_out_reg_data_35_32_sva_dfm_1_4_1_0 <= 2'b00;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_29_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= MUX_s_1_2_2((pe_manager_base_weight_sva[0]), PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      rva_out_reg_data_35_32_sva_dfm_1_4_3_2 <= rva_out_reg_data_35_32_sva_dfm_1_3[3:2];
      rva_out_reg_data_35_32_sva_dfm_1_4_1_0 <= MUX_v_2_2_2((weight_read_addrs_2_14_1_lpi_1_dfm_1[1:0]),
          (rva_out_reg_data_35_32_sva_dfm_1_3[1:0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_3 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_55_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_31_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_40_itm_1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_284_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= rva_out_reg_data_23_17_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_285_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= rva_out_reg_data_15_9_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_286_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= rva_out_reg_data_39_36_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_287_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= rva_out_reg_data_46_40_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_1_4 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_288_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_1_4 <= rva_out_reg_data_62_48_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]))) & while_stage_0_4 )
        begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_33_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_2 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_56_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ reg_rva_in_reg_rw_sva_2_cse) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= input_read_req_valid_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= 6'b000000;
      rva_out_reg_data_23_17_sva_dfm_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_175_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= MUX_v_6_2_2(6'b000000, (pe_manager_base_weight_sva_mx2[14:9]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
      rva_out_reg_data_23_17_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_base_weight_sva_mx2[7:1]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_289_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= rva_out_reg_data_15_9_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_290_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= rva_out_reg_data_35_32_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_291_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= rva_out_reg_data_39_36_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_292_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= rva_out_reg_data_46_40_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_1_3 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_293_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_1_3 <= rva_out_reg_data_62_48_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]))) & while_stage_0_4 )
        begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_182_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= rva_out_reg_data_15_9_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_294_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= rva_out_reg_data_35_32_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_295_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= rva_out_reg_data_39_36_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_296_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= rva_out_reg_data_46_40_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_48_sva_dfm_1_2 <= 15'b000000000000000;
    end
    else if ( rva_out_reg_data_and_297_enex5 ) begin
      rva_out_reg_data_62_48_sva_dfm_1_2 <= pe_manager_base_input_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (and_dcpl_488 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        & while_stage_0_3 ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_2_1,
          PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_488 & (~ (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[0]))
        & (~ (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[3]))
        & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[2])
        & and_dcpl_495 & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2))
        & (~ (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[1]))
        & and_dcpl_172 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ reg_rva_in_reg_rw_sva_st_1_1_cse) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
        & while_stage_0_3 ) begin
      input_read_req_valid_lpi_1_dfm_1_2 <= input_read_req_valid_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_1 <= 7'b0000000;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_46_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3;
      rva_out_reg_data_15_9_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_num_input_sva[7:1]),
          and_279_cse);
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_48_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_1 <= pe_config_is_cluster_sva;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= pe_config_is_bias_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (or_dcpl_121 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
        | (~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]))))
        & and_dcpl_180 ) begin
      input_read_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= 1'b0;
      rva_out_reg_data_35_32_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_39_36_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_1_1 <= 7'b0000000;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_52_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= (pe_config_num_output_sva[7]) & (~(and_279_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1))
          & PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
      rva_out_reg_data_35_32_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl
          & (signext_4_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1)) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_39_36_sva_dfm_1_1 <= (pe_manager_base_bias_sva[7:4]) & ({{3{and_279_cse}},
          and_279_cse}) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_46_40_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_6_nl
          & (signext_7_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1)) & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_15
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0
          <= 15'b000000000000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_80_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_15
          <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm[15];
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0
          <= MUX_v_15_2_2(rva_out_reg_data_62_48_sva_dfm_1_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm[14:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_0 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_170_cse ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_0 <= weight_port_read_out_data_0_1_sva_dfm_1_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_209_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_rsp_1 <= weight_port_read_out_data_0_1_sva_dfm_1_14_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_4_rsp_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_298_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_4_rsp_0 <= rva_out_reg_data_30_25_sva_dfm_3_5_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_4_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_128_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_4_rsp_1 <= rva_out_reg_data_30_25_sva_dfm_3_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_5_3_2 <= 2'b00;
      rva_out_reg_data_35_32_sva_dfm_1_5_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_150_cse ) begin
      rva_out_reg_data_35_32_sva_dfm_1_5_3_2 <= rva_out_reg_data_35_32_sva_dfm_1_4_3_2;
      rva_out_reg_data_35_32_sva_dfm_1_5_1_0 <= rva_out_reg_data_35_32_sva_dfm_1_4_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_3_5_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_299_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_3_5_2 <= rva_out_reg_data_30_25_sva_dfm_2_5_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_3_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_166_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_3_1_0 <= rva_out_reg_data_30_25_sva_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_2_5_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_300_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_2_5_2 <= rva_out_reg_data_30_25_sva_dfm_1[5:2];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_2_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_168_ssc ) begin
      rva_out_reg_data_30_25_sva_dfm_2_1_0 <= MUX_v_2_2_2((pe_manager_base_weight_sva[1:0]),
          (rva_out_reg_data_30_25_sva_dfm_1[1:0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_1_14_0 <= 15'b000000000000000;
    end
    else if ( mux_466_nl & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_0_1_sva_dfm_1_1_14_0 <= MUX1HOT_v_15_9_2(weight_port_read_out_data_0_1_sva_mx0_14_0,
          (input_mem_banks_read_read_data_lpi_1_dfm_1_4[30:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[30:16]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[30:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[30:16]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[30:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[30:16]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[30:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[14:0]),
          {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_126
          , weight_mem_run_3_for_5_and_158_ssc , weight_mem_run_3_for_5_and_159_ssc
          , weight_mem_run_3_for_5_and_160_ssc , weight_mem_run_3_for_5_and_161_ssc
          , weight_mem_run_3_for_5_and_162_cse , weight_mem_run_3_for_5_and_163_cse
          , weight_mem_run_3_for_5_and_164_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_5_rsp_0 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_164_cse ) begin
      weight_port_read_out_data_0_1_sva_dfm_5_rsp_0 <= weight_port_read_out_data_0_1_sva_dfm_4_15;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_5_rsp_1 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_210_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_5_rsp_1 <= weight_port_read_out_data_0_1_sva_dfm_4_14_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_7_rsp_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_301_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_7_rsp_0 <= rva_out_reg_data_30_25_sva_dfm_6_5_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_7_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_68_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_7_rsp_1 <= rva_out_reg_data_30_25_sva_dfm_6_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_4_15 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_166_cse ) begin
      weight_port_read_out_data_0_1_sva_dfm_4_15 <= reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_4_14_0 <= 15'b000000000000000;
    end
    else if ( weight_port_read_out_data_and_211_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_4_14_0 <= reg_weight_port_read_out_data_0_1_sva_dfm_3_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_6_5_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_302_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_6_5_2 <= reg_rva_out_reg_data_30_25_sva_dfm_5_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_6_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_89_ssc ) begin
      rva_out_reg_data_30_25_sva_dfm_6_1_0 <= reg_rva_out_reg_data_30_25_sva_dfm_5_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1_3_2 <= 2'b00;
      rva_out_reg_data_35_32_sva_dfm_4_1_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_130_ssc ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1_3_2 <= MUX1HOT_v_2_4_2(rva_out_reg_data_35_32_sva_dfm_1_5_3_2,
          rva_out_reg_data_35_32_sva_dfm_6_mx1_3_2, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[35:34]),
          (weight_port_read_out_data_0_2_sva_dfm_2[3:2]), {PECore_PushAxiRsp_if_asn_93
          , PECore_PushAxiRsp_if_asn_95 , PECore_PushAxiRsp_if_asn_91 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_35_32_sva_dfm_4_1_1_0 <= MUX1HOT_v_2_4_2(rva_out_reg_data_35_32_sva_dfm_1_5_1_0,
          rva_out_reg_data_35_32_sva_dfm_6_mx1_1_0, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[33:32]),
          (weight_port_read_out_data_0_2_sva_dfm_2[1:0]), {PECore_PushAxiRsp_if_asn_93
          , PECore_PushAxiRsp_if_asn_95 , PECore_PushAxiRsp_if_asn_91 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_6_rsp_0 <= 2'b00;
      rva_out_reg_data_35_32_sva_dfm_6_rsp_1 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_146_cse ) begin
      rva_out_reg_data_35_32_sva_dfm_6_rsp_0 <= rva_out_reg_data_35_32_sva_dfm_6_mx1_3_2;
      rva_out_reg_data_35_32_sva_dfm_6_rsp_1 <= rva_out_reg_data_35_32_sva_dfm_6_mx1_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_9_5_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_303_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_9_5_2 <= reg_rva_out_reg_data_30_25_sva_dfm_8_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_9_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_26_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_9_1_0 <= reg_rva_out_reg_data_30_25_sva_dfm_8_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_10_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_210_enex5 | rva_out_reg_data_and_191_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_10_enexo <= rva_out_reg_data_and_210_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_8_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_209_enex5 | rva_out_reg_data_and_192_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_8_enexo <= rva_out_reg_data_and_209_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_214_enex5 | rva_out_reg_data_and_193_enex5 ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_5_enexo <= rva_out_reg_data_and_214_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_215_enex5 | rva_out_reg_data_and_194_enex5 ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_5_enexo <= rva_out_reg_data_and_215_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_216_enex5 | rva_out_reg_data_and_195_enex5 ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_5_enexo <= rva_out_reg_data_and_216_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_217_enex5 | rva_out_reg_data_and_196_enex5 ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_5_enexo <= rva_out_reg_data_and_217_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_218_enex5 | rva_out_reg_data_and_197_enex5 ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_5_enexo <= rva_out_reg_data_and_218_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_219_enex5 | rva_out_reg_data_and_198_enex5 ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_5_enexo <= rva_out_reg_data_and_219_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_220_enex5 | rva_out_reg_data_and_199_enex5 ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_5_enexo <= rva_out_reg_data_and_220_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_221_enex5 | rva_out_reg_data_and_200_enex5 ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_5_enexo <= rva_out_reg_data_and_221_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_222_enex5 | rva_out_reg_data_and_201_enex5 ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_5_enexo <= rva_out_reg_data_and_222_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_223_enex5 | rva_out_reg_data_and_202_enex5 ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_5_enexo <= rva_out_reg_data_and_223_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_224_enex5 | rva_out_reg_data_and_203_enex5 ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_5_enexo <= rva_out_reg_data_and_224_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_211_enex5 | rva_out_reg_data_and_204_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_5_enexo <= rva_out_reg_data_and_211_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_225_enex5 | rva_out_reg_data_and_205_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_5_enexo <= rva_out_reg_data_and_225_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_212_enex5 | rva_out_reg_data_and_206_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_5_enexo <= rva_out_reg_data_and_212_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_213_enex5 | rva_out_reg_data_and_207_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_5_enexo <= rva_out_reg_data_and_213_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_204_enex5 | weight_port_read_out_data_and_172_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_5_enexo <= weight_port_read_out_data_and_204_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_61_enex5 | input_mem_banks_read_read_data_and_57_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_5_enexo
          <= input_mem_banks_read_read_data_and_61_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_62_enex5 | input_mem_banks_read_read_data_and_58_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_5_enexo
          <= input_mem_banks_read_read_data_and_62_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_5_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_210_enex5 | weight_port_read_out_data_and_173_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_5_1_enexo <= weight_port_read_out_data_and_210_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_63_enex5 | input_mem_banks_read_read_data_and_59_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_5_enexo
          <= input_mem_banks_read_read_data_and_63_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_64_enex5 | input_mem_banks_read_read_data_and_60_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_5_enexo
          <= input_mem_banks_read_read_data_and_64_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_vector_data_6_35_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1099_cse | accum_vector_data_and_24_enex5 ) begin
      reg_accum_vector_data_6_35_0_sva_dfm_1_1_enexo <= and_1099_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_vector_data_5_35_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1099_cse | accum_vector_data_and_25_enex5 ) begin
      reg_accum_vector_data_5_35_0_sva_dfm_1_1_enexo <= and_1099_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_vector_data_4_35_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1099_cse | accum_vector_data_and_26_enex5 ) begin
      reg_accum_vector_data_4_35_0_sva_dfm_1_1_enexo <= and_1099_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_vector_data_3_35_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1099_cse | accum_vector_data_and_27_enex5 ) begin
      reg_accum_vector_data_3_35_0_sva_dfm_1_1_enexo <= and_1099_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_vector_data_2_35_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1099_cse | accum_vector_data_and_28_enex5 ) begin
      reg_accum_vector_data_2_35_0_sva_dfm_1_1_enexo <= and_1099_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_vector_data_1_35_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1099_cse | accum_vector_data_and_29_enex5 ) begin
      reg_accum_vector_data_1_35_0_sva_dfm_1_1_enexo <= and_1099_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_vector_data_0_35_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1099_cse | accum_vector_data_and_30_enex5 ) begin
      reg_accum_vector_data_0_35_0_sva_dfm_1_1_enexo <= and_1099_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_vector_data_7_35_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1120_tmp | accum_vector_data_and_7_enex5 ) begin
      reg_accum_vector_data_7_35_0_sva_dfm_1_1_enexo <= and_1120_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_1_enex5 | input_mem_banks_read_1_read_data_and_5_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_1_read_data_and_1_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp | weight_port_read_out_data_and_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000
          <= data_in_tmp_operator_2_for_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_174_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000001
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_175_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000001
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000002
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_176_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000002
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000003
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_177_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000003
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000004
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_178_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000004
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000005
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_179_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000005
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000006
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_180_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000006
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000007
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_181_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000007
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000008
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_182_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000008
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000009
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_183_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000009
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000010
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_184_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000010
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000011
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_185_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000011
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000012
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_186_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000012
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000013
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_187_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000013
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000014
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_1_cse | weight_port_read_out_data_and_188_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000014
          <= data_in_tmp_operator_2_for_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_189_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000001
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_190_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000001
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000002
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_191_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000002
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000003
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_192_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000003
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000004
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_193_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000004
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000005
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_194_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000005
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000006
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_195_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000006
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000007
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_196_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000007
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000008
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_197_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000008
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000009
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_198_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000009
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000010
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_199_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000010
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000011
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_200_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000011
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000012
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_201_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000012
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000013
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_202_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000013
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000014
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_16_cse | weight_port_read_out_data_and_203_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_15_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000014
          <= data_in_tmp_operator_2_for_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_31_tmp | weight_port_read_out_data_and_31_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_16_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_256_255_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_3_0_16_000000
          <= data_in_tmp_operator_2_for_and_31_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_2_enex5 | input_mem_banks_read_1_read_data_and_1_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= input_mem_banks_read_1_read_data_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( weight_read_addrs_and_4_cse | weight_read_addrs_and_2_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= weight_read_addrs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= 1'b1;
    end
    else if ( weight_read_addrs_and_4_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= weight_read_addrs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3_enexo_1
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= 1'b1;
    end
    else if ( weight_read_addrs_and_4_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= weight_read_addrs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= 1'b1;
    end
    else if ( operator_15_false_1_and_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= operator_15_false_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_64_enex5 | weight_write_data_data_and_48_enex5
        ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_64_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_65_enex5 | weight_write_data_data_and_49_enex5
        ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_65_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_66_enex5 | weight_write_data_data_and_50_enex5
        ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_67_enex5 | weight_write_data_data_and_51_enex5
        ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_68_enex5 | weight_write_data_data_and_52_enex5
        ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_69_enex5 | weight_write_data_data_and_53_enex5
        ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_70_enex5 | weight_write_data_data_and_54_enex5
        ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_70_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_71_enex5 | weight_write_data_data_and_55_enex5
        ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_71_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_72_enex5 | weight_write_data_data_and_56_enex5
        ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_72_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_73_enex5 | weight_write_data_data_and_57_enex5
        ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_73_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_74_enex5 | weight_write_data_data_and_58_enex5
        ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_74_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_75_enex5 | weight_write_data_data_and_59_enex5
        ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_75_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_76_enex5 | weight_write_data_data_and_60_enex5
        ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_76_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_77_enex5 | weight_write_data_data_and_61_enex5
        ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_77_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_78_enex5 | weight_write_data_data_and_62_enex5
        ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_78_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_79_enex5 | weight_write_data_data_and_63_enex5
        ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_79_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_write_addrs_and_3_enex5 | weight_write_addrs_and_enex5 ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= weight_write_addrs_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_64_enex5 ) begin
      reg_weight_write_data_data_0_15_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_65_enex5 ) begin
      reg_weight_write_data_data_0_14_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_66_enex5 ) begin
      reg_weight_write_data_data_0_13_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_67_enex5 ) begin
      reg_weight_write_data_data_0_12_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_68_enex5 ) begin
      reg_weight_write_data_data_0_11_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_69_enex5 ) begin
      reg_weight_write_data_data_0_10_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_70_enex5 ) begin
      reg_weight_write_data_data_0_9_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_71_enex5 ) begin
      reg_weight_write_data_data_0_8_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_72_enex5 ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_73_enex5 ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_74_enex5 ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_75_enex5 ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_76_enex5 ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_77_enex5 ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_78_enex5 ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_data_data_and_79_enex5 ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_write_addrs_and_3_enex5 ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_read_addrs_and_enex5 ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_config_num_output_enexo <= 1'b1;
    end
    else if ( pe_config_num_manager_and_cse | pe_config_UpdateManagerCounter_if_if_and_enex5
        ) begin
      reg_pe_config_num_output_enexo <= pe_config_num_manager_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_16_cse | weight_read_addrs_and_27_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= while_if_and_16_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_data_sva_1_enexo <= 1'b1;
    end
    else if ( rva_in_reg_data_and_tmp | PEManager_15U_PEManagerWrite_and_enex5 )
        begin
      reg_rva_in_reg_data_sva_1_enexo <= rva_in_reg_data_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_65_enex5 | input_mem_banks_read_read_data_and_61_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_4_enexo
          <= input_mem_banks_read_read_data_and_65_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_66_enex5 | input_mem_banks_read_read_data_and_62_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_4_enexo
          <= input_mem_banks_read_read_data_and_66_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_67_enex5 | input_mem_banks_read_read_data_and_63_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_4_enexo
          <= input_mem_banks_read_read_data_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_68_enex5 | input_mem_banks_read_read_data_and_64_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_4_enexo
          <= input_mem_banks_read_read_data_and_68_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 | input_mem_banks_read_1_read_data_and_2_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_1_read_data_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_301_enex5 | rva_out_reg_data_and_208_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_7_enexo <= rva_out_reg_data_and_301_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_226_enex5 | rva_out_reg_data_and_209_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_enexo <= rva_out_reg_data_and_226_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_227_enex5 | rva_out_reg_data_and_210_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_enexo <= rva_out_reg_data_and_227_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_205_enex5 | weight_port_read_out_data_and_204_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_4_enexo <= weight_port_read_out_data_and_205_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_228_enex5 | rva_out_reg_data_and_211_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_enexo <= rva_out_reg_data_and_228_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_229_enex5 | rva_out_reg_data_and_212_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_enexo <= rva_out_reg_data_and_229_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_230_enex5 | rva_out_reg_data_and_213_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_4_enexo <= rva_out_reg_data_and_230_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_231_enex5 | rva_out_reg_data_and_214_enex5 ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_4_enexo <= rva_out_reg_data_and_231_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_232_enex5 | rva_out_reg_data_and_215_enex5 ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_4_enexo <= rva_out_reg_data_and_232_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_233_enex5 | rva_out_reg_data_and_216_enex5 ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_4_enexo <= rva_out_reg_data_and_233_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_234_enex5 | rva_out_reg_data_and_217_enex5 ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_4_enexo <= rva_out_reg_data_and_234_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_235_enex5 | rva_out_reg_data_and_218_enex5 ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_4_enexo <= rva_out_reg_data_and_235_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_236_enex5 | rva_out_reg_data_and_219_enex5 ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_4_enexo <= rva_out_reg_data_and_236_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_237_enex5 | rva_out_reg_data_and_220_enex5 ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_4_enexo <= rva_out_reg_data_and_237_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_238_enex5 | rva_out_reg_data_and_221_enex5 ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_4_enexo <= rva_out_reg_data_and_238_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_239_enex5 | rva_out_reg_data_and_222_enex5 ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_4_enexo <= rva_out_reg_data_and_239_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_240_enex5 | rva_out_reg_data_and_223_enex5 ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_4_enexo <= rva_out_reg_data_and_240_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_241_enex5 | rva_out_reg_data_and_224_enex5 ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_4_enexo <= rva_out_reg_data_and_241_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_242_enex5 | rva_out_reg_data_and_225_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_4_enexo <= rva_out_reg_data_and_242_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_69_enex5 | input_mem_banks_read_read_data_and_65_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3_enexo
          <= input_mem_banks_read_read_data_and_69_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_70_enex5 | input_mem_banks_read_read_data_and_66_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3_enexo
          <= input_mem_banks_read_read_data_and_70_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_71_enex5 | input_mem_banks_read_read_data_and_67_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3_enexo
          <= input_mem_banks_read_read_data_and_71_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_72_enex5 | input_mem_banks_read_read_data_and_68_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3_enexo
          <= input_mem_banks_read_read_data_and_72_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp | input_mem_banks_read_1_read_data_and_3_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= input_mem_banks_read_1_read_data_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_243_enex5 | rva_out_reg_data_and_226_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= rva_out_reg_data_and_243_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_244_enex5 | rva_out_reg_data_and_227_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= rva_out_reg_data_and_244_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_206_enex5 | weight_port_read_out_data_and_205_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_enexo <= weight_port_read_out_data_and_206_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_245_enex5 | rva_out_reg_data_and_228_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_3_enexo <= rva_out_reg_data_and_245_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_246_enex5 | rva_out_reg_data_and_229_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_enexo <= rva_out_reg_data_and_246_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_247_enex5 | rva_out_reg_data_and_230_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_3_enexo <= rva_out_reg_data_and_247_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_248_enex5 | rva_out_reg_data_and_231_enex5 ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_3_enexo <= rva_out_reg_data_and_248_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_249_enex5 | rva_out_reg_data_and_232_enex5 ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_3_enexo <= rva_out_reg_data_and_249_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_250_enex5 | rva_out_reg_data_and_233_enex5 ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_3_enexo <= rva_out_reg_data_and_250_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_251_enex5 | rva_out_reg_data_and_234_enex5 ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_3_enexo <= rva_out_reg_data_and_251_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_252_enex5 | rva_out_reg_data_and_235_enex5 ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_3_enexo <= rva_out_reg_data_and_252_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_253_enex5 | rva_out_reg_data_and_236_enex5 ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_3_enexo <= rva_out_reg_data_and_253_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_254_enex5 | rva_out_reg_data_and_237_enex5 ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_3_enexo <= rva_out_reg_data_and_254_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_255_enex5 | rva_out_reg_data_and_238_enex5 ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_3_enexo <= rva_out_reg_data_and_255_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_256_enex5 | rva_out_reg_data_and_239_enex5 ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_3_enexo <= rva_out_reg_data_and_256_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_257_enex5 | rva_out_reg_data_and_240_enex5 ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_3_enexo <= rva_out_reg_data_and_257_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_258_enex5 | rva_out_reg_data_and_241_enex5 ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_3_enexo <= rva_out_reg_data_and_258_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_259_enex5 | rva_out_reg_data_and_242_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_3_enexo <= rva_out_reg_data_and_259_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= 1'b1;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_1_for_and_cse | weight_mem_write_arbxbar_xbar_for_empty_and_3_enex5
        ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= weight_mem_write_arbxbar_xbar_for_1_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_73_enex5 | input_mem_banks_read_read_data_and_69_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= input_mem_banks_read_read_data_and_73_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_74_enex5 | input_mem_banks_read_read_data_and_70_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= input_mem_banks_read_read_data_and_74_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_75_enex5 | input_mem_banks_read_read_data_and_71_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= input_mem_banks_read_read_data_and_75_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_76_enex5 | input_mem_banks_read_read_data_and_72_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= input_mem_banks_read_read_data_and_76_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_261_enex5 | rva_out_reg_data_and_243_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= rva_out_reg_data_and_261_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_262_enex5 | rva_out_reg_data_and_244_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= rva_out_reg_data_and_262_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_208_enex5 | weight_port_read_out_data_and_206_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_enexo <= weight_port_read_out_data_and_208_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_209_enex5 | weight_port_read_out_data_and_207_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_209_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_263_enex5 | rva_out_reg_data_and_245_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_2_enexo <= rva_out_reg_data_and_263_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_264_enex5 | rva_out_reg_data_and_246_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_enexo <= rva_out_reg_data_and_264_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_265_enex5 | rva_out_reg_data_and_247_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_2_enexo <= rva_out_reg_data_and_265_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_266_enex5 | rva_out_reg_data_and_248_enex5 ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_2_enexo <= rva_out_reg_data_and_266_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_267_enex5 | rva_out_reg_data_and_249_enex5 ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_2_enexo <= rva_out_reg_data_and_267_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_268_enex5 | rva_out_reg_data_and_250_enex5 ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_2_enexo <= rva_out_reg_data_and_268_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_269_enex5 | rva_out_reg_data_and_251_enex5 ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_2_enexo <= rva_out_reg_data_and_269_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_270_enex5 | rva_out_reg_data_and_252_enex5 ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_2_enexo <= rva_out_reg_data_and_270_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_271_enex5 | rva_out_reg_data_and_253_enex5 ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_2_enexo <= rva_out_reg_data_and_271_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_272_enex5 | rva_out_reg_data_and_254_enex5 ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_2_enexo <= rva_out_reg_data_and_272_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_273_enex5 | rva_out_reg_data_and_255_enex5 ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_2_enexo <= rva_out_reg_data_and_273_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_274_enex5 | rva_out_reg_data_and_256_enex5 ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_2_enexo <= rva_out_reg_data_and_274_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_275_enex5 | rva_out_reg_data_and_257_enex5 ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_2_enexo <= rva_out_reg_data_and_275_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_276_enex5 | rva_out_reg_data_and_258_enex5 ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_2_enexo <= rva_out_reg_data_and_276_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_277_enex5 | rva_out_reg_data_and_259_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_2_enexo <= rva_out_reg_data_and_277_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_77_enex5 | input_mem_banks_read_read_data_and_73_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= input_mem_banks_read_read_data_and_77_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_78_enex5 | input_mem_banks_read_read_data_and_74_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo
          <= input_mem_banks_read_read_data_and_78_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_79_enex5 | input_mem_banks_read_read_data_and_75_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= input_mem_banks_read_read_data_and_79_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_80_enex5 | input_mem_banks_read_read_data_and_76_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= input_mem_banks_read_read_data_and_80_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_298_enex5 | rva_out_reg_data_and_260_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_4_enexo <= rva_out_reg_data_and_298_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_278_enex5 | rva_out_reg_data_and_261_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_4_enexo <= rva_out_reg_data_and_278_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_279_enex5 | rva_out_reg_data_and_262_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_6_enexo <= rva_out_reg_data_and_279_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_127_tmp | weight_port_read_out_data_and_208_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_1_enexo <= weight_port_read_out_data_and_127_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1344_cse | rva_out_reg_data_and_263_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_4_1_enexo <= and_1344_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1344_cse | rva_out_reg_data_and_264_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_enexo <= and_1344_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1344_cse | rva_out_reg_data_and_265_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_4_1_enexo <= and_1344_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_266_enex5 ) begin
      reg_rva_out_reg_data_255_240_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_267_enex5 ) begin
      reg_rva_out_reg_data_239_224_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_268_enex5 ) begin
      reg_rva_out_reg_data_223_208_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_269_enex5 ) begin
      reg_rva_out_reg_data_207_192_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_270_enex5 ) begin
      reg_rva_out_reg_data_191_176_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_271_enex5 ) begin
      reg_rva_out_reg_data_175_160_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_272_enex5 ) begin
      reg_rva_out_reg_data_159_144_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_273_enex5 ) begin
      reg_rva_out_reg_data_143_128_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_274_enex5 ) begin
      reg_rva_out_reg_data_127_112_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_275_enex5 ) begin
      reg_rva_out_reg_data_111_96_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_276_enex5 ) begin
      reg_rva_out_reg_data_95_80_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_cse | rva_out_reg_data_and_277_enex5 ) begin
      reg_rva_out_reg_data_79_64_sva_dfm_4_1_enexo <= rva_out_reg_data_and_134_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_54_tmp | input_mem_banks_read_read_data_and_77_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_read_data_and_54_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_54_tmp | input_mem_banks_read_read_data_and_78_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_1 <= input_mem_banks_read_read_data_and_54_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_54_tmp | input_mem_banks_read_read_data_and_79_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_2 <= input_mem_banks_read_read_data_and_54_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_3 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_54_tmp | input_mem_banks_read_read_data_and_80_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo_3 <= input_mem_banks_read_read_data_and_54_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_282_enex5 | rva_out_reg_data_and_278_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_3_enexo <= rva_out_reg_data_and_282_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_283_enex5 | rva_out_reg_data_and_279_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_5_enexo <= rva_out_reg_data_and_283_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_287_enex5 | rva_out_reg_data_and_280_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_4_enexo <= rva_out_reg_data_and_287_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_286_enex5 | rva_out_reg_data_and_281_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_4_enexo <= rva_out_reg_data_and_286_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_284_enex5 | rva_out_reg_data_and_282_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_2_enexo <= rva_out_reg_data_and_284_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_285_enex5 | rva_out_reg_data_and_283_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_4_enexo <= rva_out_reg_data_and_285_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_56_enex5 | input_mem_banks_read_read_data_and_55_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_read_data_and_56_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_175_cse | rva_out_reg_data_and_284_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= rva_out_reg_data_and_175_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_289_enex5 | rva_out_reg_data_and_285_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= rva_out_reg_data_and_289_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_291_enex5 | rva_out_reg_data_and_286_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= rva_out_reg_data_and_291_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_292_enex5 | rva_out_reg_data_and_287_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= rva_out_reg_data_and_292_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_293_enex5 | rva_out_reg_data_and_288_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_1_3_enexo <= rva_out_reg_data_and_293_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_tmp | input_mem_banks_read_read_data_and_56_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo_1 <= input_mem_banks_read_1_read_data_and_4_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_182_enex5 | rva_out_reg_data_and_289_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= rva_out_reg_data_and_182_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_294_enex5 | rva_out_reg_data_and_290_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= rva_out_reg_data_and_294_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_295_enex5 | rva_out_reg_data_and_291_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= rva_out_reg_data_and_295_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_296_enex5 | rva_out_reg_data_and_292_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= rva_out_reg_data_and_296_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_297_enex5 | rva_out_reg_data_and_293_enex5 ) begin
      reg_rva_out_reg_data_62_48_sva_dfm_1_2_enexo <= rva_out_reg_data_and_297_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_46_cse | rva_out_reg_data_and_182_enex5
        ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_46_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_52_cse | rva_out_reg_data_and_294_enex5
        ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_52_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_52_cse | rva_out_reg_data_and_295_enex5
        ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_52_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_52_cse | rva_out_reg_data_and_296_enex5
        ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_52_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_input_enexo <= 1'b1;
    end
    else if ( pe_manager_base_input_and_tmp | rva_out_reg_data_and_297_enex5 ) begin
      reg_pe_manager_base_input_enexo <= pe_manager_base_input_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1266_cse | weight_port_read_out_data_and_209_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_1_enexo <= and_1266_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_299_enex5 | rva_out_reg_data_and_298_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_3_enexo <= rva_out_reg_data_and_299_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_300_enex5 | rva_out_reg_data_and_299_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_2_enexo <= rva_out_reg_data_and_300_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_175_cse | rva_out_reg_data_and_300_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= rva_out_reg_data_and_175_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_211_enex5 | weight_port_read_out_data_and_210_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_4_1_enexo <= weight_port_read_out_data_and_211_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_302_enex5 | rva_out_reg_data_and_301_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= rva_out_reg_data_and_302_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_207_enex5 | weight_port_read_out_data_and_211_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_207_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_260_enex5 | rva_out_reg_data_and_302_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= rva_out_reg_data_and_260_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_8_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_208_enex5 | rva_out_reg_data_and_303_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_8_enexo <= rva_out_reg_data_and_208_enex5;
    end
  end
  assign nl_operator_4_false_acc_nl = pe_config_manager_counter_sva_mx1 + 4'b0001;
  assign operator_4_false_acc_nl = nl_operator_4_false_acc_nl[3:0];
  assign pe_config_UpdateManagerCounter_if_not_7_nl = ~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  assign nl_input_read_addrs_sva_1_1  = pe_config_input_counter_sva_mx1 + (pe_manager_base_input_sva_mx1[7:0]);
  assign PECore_UpdateFSM_switch_lp_not_25_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_11;
  assign PECore_UpdateFSM_switch_lp_not_26_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_11;
  assign PECore_UpdateFSM_switch_lp_not_27_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_11;
  assign PECore_UpdateFSM_switch_lp_not_28_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_11;
  assign PECore_UpdateFSM_switch_lp_not_29_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_11;
  assign PECore_UpdateFSM_switch_lp_not_30_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_11;
  assign PECore_UpdateFSM_switch_lp_not_19_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_11;
  assign nl_ProductSum_for_acc_41_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_24_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_23_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_22_z);
  assign ProductSum_for_acc_41_nl = nl_ProductSum_for_acc_41_nl[35:0];
  assign nl_ProductSum_for_acc_42_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_21_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_20_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_19_z);
  assign ProductSum_for_acc_42_nl = nl_ProductSum_for_acc_42_nl[35:0];
  assign nl_ProductSum_for_acc_43_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_18_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_17_z);
  assign ProductSum_for_acc_43_nl = nl_ProductSum_for_acc_43_nl[34:0];
  assign nl_ProductSum_for_acc_40_nl = ProductSum_for_acc_41_nl + ProductSum_for_acc_42_nl
      + conv_u2s_35_36(ProductSum_for_acc_43_nl);
  assign ProductSum_for_acc_40_nl = nl_ProductSum_for_acc_40_nl[35:0];
  assign PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_nl = MUX_v_36_2_2(accum_vector_data_6_35_0_sva,
      ProductSum_for_acc_40_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_9);
  assign PECore_UpdateFSM_switch_lp_not_31_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_33_nl = conv_u2u_34_36(Datapath_for_6_ProductSum_for_acc_1_1)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_39_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_38_z);
  assign ProductSum_for_acc_33_nl = nl_ProductSum_for_acc_33_nl[35:0];
  assign nl_ProductSum_for_acc_34_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_37_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_36_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_35_z);
  assign ProductSum_for_acc_34_nl = nl_ProductSum_for_acc_34_nl[35:0];
  assign nl_ProductSum_for_acc_35_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_34_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_33_z);
  assign ProductSum_for_acc_35_nl = nl_ProductSum_for_acc_35_nl[34:0];
  assign nl_ProductSum_for_acc_32_nl = ProductSum_for_acc_33_nl + ProductSum_for_acc_34_nl
      + conv_u2s_35_36(ProductSum_for_acc_35_nl);
  assign ProductSum_for_acc_32_nl = nl_ProductSum_for_acc_32_nl[35:0];
  assign PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_1_nl = MUX_v_36_2_2(accum_vector_data_5_35_0_sva,
      ProductSum_for_acc_32_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_9);
  assign PECore_UpdateFSM_switch_lp_not_32_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_25_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_56_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_55_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_54_z);
  assign ProductSum_for_acc_25_nl = nl_ProductSum_for_acc_25_nl[35:0];
  assign nl_ProductSum_for_acc_26_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_53_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_52_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_51_z);
  assign ProductSum_for_acc_26_nl = nl_ProductSum_for_acc_26_nl[35:0];
  assign nl_ProductSum_for_acc_27_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_50_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_49_z);
  assign ProductSum_for_acc_27_nl = nl_ProductSum_for_acc_27_nl[34:0];
  assign nl_ProductSum_for_acc_24_nl = ProductSum_for_acc_25_nl + ProductSum_for_acc_26_nl
      + conv_u2s_35_36(ProductSum_for_acc_27_nl);
  assign ProductSum_for_acc_24_nl = nl_ProductSum_for_acc_24_nl[35:0];
  assign PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_2_nl = MUX_v_36_2_2(accum_vector_data_4_35_0_sva,
      ProductSum_for_acc_24_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_9);
  assign PECore_UpdateFSM_switch_lp_not_33_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_21_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_63_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_62_z);
  assign ProductSum_for_acc_21_nl = nl_ProductSum_for_acc_21_nl[35:0];
  assign nl_ProductSum_for_acc_22_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_61_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_60_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_59_z);
  assign ProductSum_for_acc_22_nl = nl_ProductSum_for_acc_22_nl[35:0];
  assign nl_ProductSum_for_acc_23_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_58_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_57_z);
  assign ProductSum_for_acc_23_nl = nl_ProductSum_for_acc_23_nl[34:0];
  assign nl_ProductSum_for_acc_20_nl = ProductSum_for_acc_21_nl + ProductSum_for_acc_22_nl
      + conv_u2s_35_36(ProductSum_for_acc_23_nl);
  assign ProductSum_for_acc_20_nl = nl_ProductSum_for_acc_20_nl[35:0];
  assign PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_3_nl = MUX_v_36_2_2(accum_vector_data_3_35_0_sva,
      ProductSum_for_acc_20_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_9);
  assign PECore_UpdateFSM_switch_lp_not_34_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_29_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_48_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_47_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_46_z);
  assign ProductSum_for_acc_29_nl = nl_ProductSum_for_acc_29_nl[35:0];
  assign nl_ProductSum_for_acc_30_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_45_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_44_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_43_z);
  assign ProductSum_for_acc_30_nl = nl_ProductSum_for_acc_30_nl[35:0];
  assign nl_ProductSum_for_acc_31_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_42_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_41_z);
  assign ProductSum_for_acc_31_nl = nl_ProductSum_for_acc_31_nl[34:0];
  assign nl_ProductSum_for_acc_28_nl = ProductSum_for_acc_29_nl + ProductSum_for_acc_30_nl
      + conv_u2s_35_36(ProductSum_for_acc_31_nl);
  assign ProductSum_for_acc_28_nl = nl_ProductSum_for_acc_28_nl[35:0];
  assign PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_4_nl = MUX_v_36_2_2(accum_vector_data_2_35_0_sva,
      ProductSum_for_acc_28_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_9);
  assign PECore_UpdateFSM_switch_lp_not_35_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_37_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_32_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_31_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_30_z);
  assign ProductSum_for_acc_37_nl = nl_ProductSum_for_acc_37_nl[35:0];
  assign nl_ProductSum_for_acc_38_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_29_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_28_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_27_z);
  assign ProductSum_for_acc_38_nl = nl_ProductSum_for_acc_38_nl[35:0];
  assign nl_ProductSum_for_acc_39_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_26_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_25_z);
  assign ProductSum_for_acc_39_nl = nl_ProductSum_for_acc_39_nl[34:0];
  assign nl_ProductSum_for_acc_36_nl = ProductSum_for_acc_37_nl + ProductSum_for_acc_38_nl
      + conv_u2s_35_36(ProductSum_for_acc_39_nl);
  assign ProductSum_for_acc_36_nl = nl_ProductSum_for_acc_36_nl[35:0];
  assign PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_5_nl = MUX_v_36_2_2(accum_vector_data_1_35_0_sva,
      ProductSum_for_acc_36_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_9);
  assign PECore_UpdateFSM_switch_lp_not_36_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_45_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_16_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_15_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_14_z);
  assign ProductSum_for_acc_45_nl = nl_ProductSum_for_acc_45_nl[35:0];
  assign nl_ProductSum_for_acc_46_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_13_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_12_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_11_z);
  assign ProductSum_for_acc_46_nl = nl_ProductSum_for_acc_46_nl[35:0];
  assign nl_ProductSum_for_acc_47_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_10_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_9_z);
  assign ProductSum_for_acc_47_nl = nl_ProductSum_for_acc_47_nl[34:0];
  assign nl_ProductSum_for_acc_44_nl = ProductSum_for_acc_45_nl + ProductSum_for_acc_46_nl
      + conv_u2s_35_36(ProductSum_for_acc_47_nl);
  assign ProductSum_for_acc_44_nl = nl_ProductSum_for_acc_44_nl[35:0];
  assign PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_6_nl = MUX_v_36_2_2(accum_vector_data_0_35_0_sva,
      ProductSum_for_acc_44_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_9);
  assign PECore_UpdateFSM_switch_lp_not_21_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign nl_ProductSum_for_acc_48_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_8_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_7_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_6_z);
  assign ProductSum_for_acc_48_nl = nl_ProductSum_for_acc_48_nl[35:0];
  assign nl_ProductSum_for_acc_49_nl = conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_5_z)
      + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_4_z) + conv_u2u_34_36(Datapath_for_4_ProductSum_for_acc_9_cmp_3_z);
  assign ProductSum_for_acc_49_nl = nl_ProductSum_for_acc_49_nl[35:0];
  assign nl_ProductSum_for_acc_50_nl = conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_2_z)
      + conv_u2u_34_35(Datapath_for_4_ProductSum_for_acc_9_cmp_1_z);
  assign ProductSum_for_acc_50_nl = nl_ProductSum_for_acc_50_nl[34:0];
  assign nl_ProductSum_for_acc_nl = ProductSum_for_acc_48_nl + ProductSum_for_acc_49_nl
      + conv_u2s_35_36(ProductSum_for_acc_50_nl);
  assign ProductSum_for_acc_nl = nl_ProductSum_for_acc_nl[35:0];
  assign PECore_RunMac_PECore_RunMac_PECore_RunMac_mux_7_nl = MUX_v_36_2_2(accum_vector_data_7_35_0_sva,
      ProductSum_for_acc_nl, PECore_RunMac_PECore_RunMac_if_and_svs_st_8);
  assign PECore_UpdateFSM_switch_lp_not_10_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign weight_mem_run_3_for_5_and_166_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_167_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_168_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_169_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_170_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_172_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign or_1188_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_110_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_111_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_112_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_113_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_116_itm_2;
  assign mux_354_nl = MUX_s_1_2_2(or_1189_cse, or_1188_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign weight_mem_run_3_for_5_and_174_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_175_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_176_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_104_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_177_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_179_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_180_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign or_1190_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_102_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_103_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_104_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_105_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_107_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_108_itm_2;
  assign mux_355_nl = MUX_s_1_2_2(or_1189_cse, or_1190_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_nl = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[255:240]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[255:240]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[239:224]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_369
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_1_nl = MUX1HOT_v_16_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[255:240]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[255:240]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[255:240]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[255:240]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_255_16_mx0[239:224]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_371
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_130_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_131_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_252_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_133_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_254_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_255_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1});
  assign nor_510_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ or_tmp_441));
  assign mux_376_nl = MUX_s_1_2_2(nor_510_nl, or_tmp_441, or_1284_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_48_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[15:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl);
  assign and_64_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1));
  assign mux_4_nl = MUX_s_1_2_2(and_64_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_766_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_127_itm_1;
  assign or_13_nl = (~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign mux_5_nl = MUX_s_1_2_2(mux_4_nl, and_766_nl, or_13_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_138_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_80_nl
      = MUX_v_16_2_2(16'b0000000000000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[15:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_138_nl);
  assign nor_328_nl = ~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_6_nl = MUX_s_1_2_2(nor_328_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_118_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_7_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_3, (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_80_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign nor_511_nl = ~((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign nor_512_nl = ~((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | (~ reg_rva_in_reg_rw_sva_st_1_1_cse));
  assign mux_377_nl = MUX_s_1_2_2(nor_511_nl, nor_512_nl, while_stage_0_3);
  assign mux_378_nl = MUX_s_1_2_2(mux_377_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2,
      while_stage_0_4);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl
      = MUX_v_11_2_2(11'b00000000000, PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl
      = MUX_v_4_2_2(4'b0000, pe_config_manager_counter_sva_mx1, PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign and_622_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & and_dcpl_183 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]));
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl = (state_mux_1_cse!=2'b00)
      | state_0_sva_mx1;
  assign PECore_UpdateFSM_switch_lp_or_nl = PECore_UpdateFSM_switch_lp_equal_tmp_6
      | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  assign PECore_UpdateFSM_switch_lp_mux1h_16_nl = MUX1HOT_v_2_3_2((signext_2_1(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl)),
      2'b01, 2'b10, {PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      , PECore_UpdateFSM_switch_lp_or_nl , PECore_RunScale_PECore_RunScale_if_and_1_svs_1});
  assign PECore_UpdateFSM_switch_lp_nor_8_nl = ~(PECore_PushOutput_PECore_PushOutput_if_and_svs_1
      | PECore_UpdateFSM_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_and_1_nl = MUX_v_2_2_2(2'b00, PECore_UpdateFSM_switch_lp_mux1h_16_nl,
      PECore_UpdateFSM_switch_lp_nor_8_nl);
  assign mux_379_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_3_1, nor_523_cse,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_380_nl = MUX_s_1_2_2(and_1437_cse, nor_523_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nl_operator_8_false_acc_sdt_sva_1  = conv_u2s_8_9(pe_config_num_output_sva)
      + 9'b111111111;
  assign PECore_UpdateFSM_switch_lp_not_11_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign nor_525_nl = ~(PECore_RunMac_PECore_RunMac_if_and_svs_st_10 | (~(PECore_RunScale_PECore_RunScale_if_and_1_svs_10
      & mux_tmp_376)));
  assign mux_390_nl = MUX_s_1_2_2(nor_525_nl, mux_tmp_376, PECore_UpdateFSM_switch_lp_equal_tmp_2_10);
  assign mux1h_7_nl = MUX1HOT_v_15_7_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_14_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1[14:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1[14:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1[14:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[30:16]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[30:16]),
      weight_port_read_out_data_0_1_sva_mx0_14_0, {and_1017_cse , and_1018_cse ,
      and_1019_cse , and_1020_cse , and_1021_cse , and_1022_cse , nor_472_cse});
  assign not_2496_nl = ~ or_dcpl;
  assign or_1326_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1;
  assign or_1325_nl = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1;
  assign mux_394_nl = MUX_s_1_2_2(or_1326_nl, or_1325_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign or_1324_nl = nor_526_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_256_itm_1;
  assign mux_395_nl = MUX_s_1_2_2(mux_394_nl, or_1324_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]);
  assign mux_396_nl = MUX_s_1_2_2(nand_72_cse, mux_395_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign mux_36_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_3_lpi_1_dfm_1, (~ or_tmp_35),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_1335_nl = reg_weight_mem_run_3_for_5_and_146_itm_2_cse | reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_148_itm_2_cse | reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      | weight_mem_run_3_for_5_and_150_itm_2 | weight_mem_run_3_for_5_and_151_itm_2
      | reg_weight_mem_run_3_for_5_and_152_itm_2_cse | and_1441_cse;
  assign and_1442_nl = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign and_1443_nl = ((~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign mux_397_nl = MUX_s_1_2_2(and_1442_nl, and_1443_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign and_1444_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_26_itm_1)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign mux_398_nl = MUX_s_1_2_2(mux_397_nl, and_1444_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_1333_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_212_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_231_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_126_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_itm_1 | mux_398_nl;
  assign mux_399_nl = MUX_s_1_2_2(or_1335_nl, or_1333_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_260_nl = (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  assign mux_37_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_6_lpi_1_dfm_1, (~ rva_in_reg_rw_sva_st_1_4),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_136_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_215_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_18_nl
      = ~((weight_read_addrs_3_lpi_1_dfm_2_2_0!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_204_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_190_nl = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_28_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign or_189_nl = PECore_RunMac_PECore_RunMac_if_and_svs_st_2 | (~(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1
      | Arbiter_8U_Roundrobin_pick_1_if_1_and_30_tmp)) | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign mux_40_nl = MUX_s_1_2_2(or_189_nl, or_188_cse, Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp);
  assign or_182_nl = (~(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse))
      | (~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign or_180_nl = Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp;
  assign mux_38_nl = MUX_s_1_2_2(or_182_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3,
      or_180_nl);
  assign mux_41_nl = MUX_s_1_2_2(mux_40_nl, mux_38_nl, while_stage_0_5);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl
      = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]), pe_config_is_zero_first_sva_mx1,
      PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_27_nl
      = MUX_s_1_2_2(PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl,
      pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_or_5_cse_1);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_234_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_249_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_174_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_189_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_204_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_219_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_235_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_250_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_175_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_190_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_205_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_220_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_236_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_251_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_176_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_191_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_206_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_221_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_237_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_252_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_177_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_192_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_207_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_222_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_238_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_253_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_178_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_193_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_208_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_223_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_239_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_254_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_179_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_194_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_209_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_224_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_240_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_255_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_180_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_195_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_210_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_225_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_241_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_256_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_181_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_196_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_211_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_226_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_242_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_257_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_182_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_197_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_212_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_227_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_243_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_258_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_183_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_198_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_213_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_228_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_244_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_259_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_184_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_199_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_214_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_229_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_245_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_260_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_185_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_200_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_215_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_230_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_246_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_247_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign mux1h_2_nl = MUX1HOT_v_16_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[63:48]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[63:48]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[63:48]),
      {and_1025_cse , and_1026_cse , and_1027_cse});
  assign not_2436_nl = ~ or_dcpl_719;
  assign mux1h_3_nl = MUX1HOT_v_16_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[47:32]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[47:32]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[47:32]),
      {and_1025_cse , and_1026_cse , and_1027_cse});
  assign not_2438_nl = ~ or_dcpl_719;
  assign mux1h_4_nl = MUX1HOT_v_16_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[31:16]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[31:16]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[31:16]),
      {and_1025_cse , and_1026_cse , and_1027_cse});
  assign not_2440_nl = ~ or_dcpl_719;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_201_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_202_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_203_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_231_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_233_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_232_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_140_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign and_669_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign and_670_nl = and_dcpl_657 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign and_672_nl = (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      & weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_675_nl = and_dcpl_664 & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1));
  assign and_678_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_load_store_for_else_mux1h_89_nl = MUX1HOT_v_16_5_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[15:0]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[15:0]), (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[15:0]),
      (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[15:0]), (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[15:0]),
      {and_669_nl , and_670_nl , and_672_nl , and_675_nl , and_678_nl});
  assign and_668_nl = nor_335_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign weight_mem_banks_load_store_for_else_or_nl = MUX_v_16_2_2(weight_mem_banks_load_store_for_else_mux1h_89_nl,
      16'b1111111111111111, and_668_nl);
  assign and_1061_nl = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & and_dcpl_664;
  assign nor_471_nl = ~((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]) | (~ nor_335_cse));
  assign mux_340_nl = MUX_s_1_2_2(and_1061_nl, nor_471_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_348_nl = MUX_v_16_2_2(weight_mem_banks_load_store_for_else_or_nl, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[15:0]),
      mux_340_nl);
  assign nand_67_nl = ~(or_dcpl_719 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_206_nl = (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign mux_48_nl = MUX_s_1_2_2(or_206_nl, mux_tmp_46, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_205_nl = (~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign mux_47_nl = MUX_s_1_2_2(or_205_nl, mux_tmp_46, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_200_nl = (~((~(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign mux_49_nl = MUX_s_1_2_2(mux_48_nl, mux_47_nl, or_200_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_135_nl = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_134_nl = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b110)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_132_nl = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b011)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b101)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_114_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_359_itm_1
      & (pe_manager_base_weight_sva[1:0]==2'b01) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign mux_50_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, (~ pe_manager_base_weight_slc_pe_manager_base_weight_2_0_363_itm_1),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign nor_339_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | mux_tmp_51);
  assign mux_52_nl = MUX_s_1_2_2(or_tmp_59, nor_339_nl, weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1);
  assign mux_53_nl = MUX_s_1_2_2(mux_52_nl, or_tmp_59, weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign and_1062_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & fsm_output;
  assign input_mem_banks_read_1_for_mux_nl = MUX_v_8_2_2(input_read_addrs_sva_1_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4,
      and_1062_nl);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_17_nl
      = pe_manager_base_input_sva_mx1 & ({{14{and_279_cse}}, and_279_cse}) & ({{14{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
  assign or_834_nl = or_dcpl_129 | or_dcpl_700;
  assign or_160_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  assign mux_54_nl = MUX_s_1_2_2(and_dcpl_321, or_160_nl, weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]);
  assign weight_port_read_out_data_mux_67_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_26_mx0w2,
      (weight_port_read_out_data_0_3_sva_dfm_2[15]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign mux1h_1_nl = MUX1HOT_s_1_7_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_itm_1_15,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_17_itm_1[15]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_49_itm_1[15]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_81_itm_1[15]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[31]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[31]),
      weight_port_read_out_data_0_1_sva_mx0_15, {and_1017_cse , and_1018_cse , and_1019_cse
      , and_1020_cse , and_1021_cse , and_1022_cse , nor_472_cse});
  assign and_688_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign nor_463_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_3_itm_2,
      pe_manager_base_weight_sva_mx3_0, PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2,
      (pe_manager_base_weight_sva_mx2[8]), PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl =
      (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl = MUX_s_1_2_2(pe_config_is_valid_sva,
      pe_manager_zero_active_sva, and_279_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl = MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1,
      (pe_manager_num_input_sva[0]), and_279_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_1_nl = MUX_v_4_2_2(pe_config_num_manager_sva,
      (pe_manager_base_bias_sva[3:0]), and_279_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_6_nl = MUX_v_7_2_2((pe_config_num_output_sva[6:0]),
      (pe_manager_base_bias_sva[14:8]), and_279_cse);
  assign or_1448_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_14_itm_2
      | reg_weight_mem_run_3_for_5_and_146_itm_2_cse | reg_weight_mem_run_3_for_5_and_147_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_148_itm_2_cse | reg_weight_mem_run_3_for_5_and_149_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_122_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_123_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_124_itm_2;
  assign mux_466_nl = MUX_s_1_2_2(or_1189_cse, or_1448_nl, weight_mem_run_3_for_land_1_lpi_1_dfm_3);

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_9_2;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [8:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_8_2;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [7:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    result = result | (input_5 & {11{sel[5]}});
    result = result | (input_6 & {11{sel[6]}});
    result = result | (input_7 & {11{sel[7]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_3_2;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [2:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | (input_1 & {15{sel[1]}});
    result = result | (input_2 & {15{sel[2]}});
    MUX1HOT_v_15_3_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_4_2;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [3:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | (input_1 & {15{sel[1]}});
    result = result | (input_2 & {15{sel[2]}});
    result = result | (input_3 & {15{sel[3]}});
    MUX1HOT_v_15_4_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_7_2;
    input [14:0] input_6;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [6:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | (input_1 & {15{sel[1]}});
    result = result | (input_2 & {15{sel[2]}});
    result = result | (input_3 & {15{sel[3]}});
    result = result | (input_4 & {15{sel[4]}});
    result = result | (input_5 & {15{sel[5]}});
    result = result | (input_6 & {15{sel[6]}});
    MUX1HOT_v_15_7_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_9_2;
    input [14:0] input_8;
    input [14:0] input_7;
    input [14:0] input_6;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [8:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | (input_1 & {15{sel[1]}});
    result = result | (input_2 & {15{sel[2]}});
    result = result | (input_3 & {15{sel[3]}});
    result = result | (input_4 & {15{sel[4]}});
    result = result | (input_5 & {15{sel[5]}});
    result = result | (input_6 & {15{sel[6]}});
    result = result | (input_7 & {15{sel[7]}});
    result = result | (input_8 & {15{sel[8]}});
    MUX1HOT_v_15_9_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_5_2;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [4:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    MUX1HOT_v_16_5_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_6_2;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [5:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    MUX1HOT_v_16_6_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_7_2;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [6:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    MUX1HOT_v_16_7_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_8_2;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [7:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    result = result | (input_7 & {16{sel[7]}});
    MUX1HOT_v_16_8_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_9_2;
    input [15:0] input_8;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [8:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    result = result | (input_7 & {16{sel[7]}});
    result = result | (input_8 & {16{sel[8]}});
    MUX1HOT_v_16_9_2 = result;
  end
  endfunction


  function automatic [255:0] MUX1HOT_v_256_3_2;
    input [255:0] input_2;
    input [255:0] input_1;
    input [255:0] input_0;
    input [2:0] sel;
    reg [255:0] result;
  begin
    result = input_0 & {256{sel[0]}};
    result = result | (input_1 & {256{sel[1]}});
    result = result | (input_2 & {256{sel[2]}});
    MUX1HOT_v_256_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | (input_1 & {32{sel[1]}});
    result = result | (input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_8_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input [2:0] sel;
    reg  result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_s_1_8_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_8_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [10:0] input_2;
    input [10:0] input_3;
    input [10:0] input_4;
    input [10:0] input_5;
    input [10:0] input_6;
    input [10:0] input_7;
    input [2:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_11_8_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input  sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input  sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_8_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [2:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_16_8_2 = result;
  end
  endfunction


  function automatic [239:0] MUX_v_240_2_2;
    input [239:0] input_0;
    input [239:0] input_1;
    input  sel;
    reg [239:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_240_2_2 = result;
  end
  endfunction


  function automatic [255:0] MUX_v_256_256_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [255:0] input_2;
    input [255:0] input_3;
    input [255:0] input_4;
    input [255:0] input_5;
    input [255:0] input_6;
    input [255:0] input_7;
    input [255:0] input_8;
    input [255:0] input_9;
    input [255:0] input_10;
    input [255:0] input_11;
    input [255:0] input_12;
    input [255:0] input_13;
    input [255:0] input_14;
    input [255:0] input_15;
    input [255:0] input_16;
    input [255:0] input_17;
    input [255:0] input_18;
    input [255:0] input_19;
    input [255:0] input_20;
    input [255:0] input_21;
    input [255:0] input_22;
    input [255:0] input_23;
    input [255:0] input_24;
    input [255:0] input_25;
    input [255:0] input_26;
    input [255:0] input_27;
    input [255:0] input_28;
    input [255:0] input_29;
    input [255:0] input_30;
    input [255:0] input_31;
    input [255:0] input_32;
    input [255:0] input_33;
    input [255:0] input_34;
    input [255:0] input_35;
    input [255:0] input_36;
    input [255:0] input_37;
    input [255:0] input_38;
    input [255:0] input_39;
    input [255:0] input_40;
    input [255:0] input_41;
    input [255:0] input_42;
    input [255:0] input_43;
    input [255:0] input_44;
    input [255:0] input_45;
    input [255:0] input_46;
    input [255:0] input_47;
    input [255:0] input_48;
    input [255:0] input_49;
    input [255:0] input_50;
    input [255:0] input_51;
    input [255:0] input_52;
    input [255:0] input_53;
    input [255:0] input_54;
    input [255:0] input_55;
    input [255:0] input_56;
    input [255:0] input_57;
    input [255:0] input_58;
    input [255:0] input_59;
    input [255:0] input_60;
    input [255:0] input_61;
    input [255:0] input_62;
    input [255:0] input_63;
    input [255:0] input_64;
    input [255:0] input_65;
    input [255:0] input_66;
    input [255:0] input_67;
    input [255:0] input_68;
    input [255:0] input_69;
    input [255:0] input_70;
    input [255:0] input_71;
    input [255:0] input_72;
    input [255:0] input_73;
    input [255:0] input_74;
    input [255:0] input_75;
    input [255:0] input_76;
    input [255:0] input_77;
    input [255:0] input_78;
    input [255:0] input_79;
    input [255:0] input_80;
    input [255:0] input_81;
    input [255:0] input_82;
    input [255:0] input_83;
    input [255:0] input_84;
    input [255:0] input_85;
    input [255:0] input_86;
    input [255:0] input_87;
    input [255:0] input_88;
    input [255:0] input_89;
    input [255:0] input_90;
    input [255:0] input_91;
    input [255:0] input_92;
    input [255:0] input_93;
    input [255:0] input_94;
    input [255:0] input_95;
    input [255:0] input_96;
    input [255:0] input_97;
    input [255:0] input_98;
    input [255:0] input_99;
    input [255:0] input_100;
    input [255:0] input_101;
    input [255:0] input_102;
    input [255:0] input_103;
    input [255:0] input_104;
    input [255:0] input_105;
    input [255:0] input_106;
    input [255:0] input_107;
    input [255:0] input_108;
    input [255:0] input_109;
    input [255:0] input_110;
    input [255:0] input_111;
    input [255:0] input_112;
    input [255:0] input_113;
    input [255:0] input_114;
    input [255:0] input_115;
    input [255:0] input_116;
    input [255:0] input_117;
    input [255:0] input_118;
    input [255:0] input_119;
    input [255:0] input_120;
    input [255:0] input_121;
    input [255:0] input_122;
    input [255:0] input_123;
    input [255:0] input_124;
    input [255:0] input_125;
    input [255:0] input_126;
    input [255:0] input_127;
    input [255:0] input_128;
    input [255:0] input_129;
    input [255:0] input_130;
    input [255:0] input_131;
    input [255:0] input_132;
    input [255:0] input_133;
    input [255:0] input_134;
    input [255:0] input_135;
    input [255:0] input_136;
    input [255:0] input_137;
    input [255:0] input_138;
    input [255:0] input_139;
    input [255:0] input_140;
    input [255:0] input_141;
    input [255:0] input_142;
    input [255:0] input_143;
    input [255:0] input_144;
    input [255:0] input_145;
    input [255:0] input_146;
    input [255:0] input_147;
    input [255:0] input_148;
    input [255:0] input_149;
    input [255:0] input_150;
    input [255:0] input_151;
    input [255:0] input_152;
    input [255:0] input_153;
    input [255:0] input_154;
    input [255:0] input_155;
    input [255:0] input_156;
    input [255:0] input_157;
    input [255:0] input_158;
    input [255:0] input_159;
    input [255:0] input_160;
    input [255:0] input_161;
    input [255:0] input_162;
    input [255:0] input_163;
    input [255:0] input_164;
    input [255:0] input_165;
    input [255:0] input_166;
    input [255:0] input_167;
    input [255:0] input_168;
    input [255:0] input_169;
    input [255:0] input_170;
    input [255:0] input_171;
    input [255:0] input_172;
    input [255:0] input_173;
    input [255:0] input_174;
    input [255:0] input_175;
    input [255:0] input_176;
    input [255:0] input_177;
    input [255:0] input_178;
    input [255:0] input_179;
    input [255:0] input_180;
    input [255:0] input_181;
    input [255:0] input_182;
    input [255:0] input_183;
    input [255:0] input_184;
    input [255:0] input_185;
    input [255:0] input_186;
    input [255:0] input_187;
    input [255:0] input_188;
    input [255:0] input_189;
    input [255:0] input_190;
    input [255:0] input_191;
    input [255:0] input_192;
    input [255:0] input_193;
    input [255:0] input_194;
    input [255:0] input_195;
    input [255:0] input_196;
    input [255:0] input_197;
    input [255:0] input_198;
    input [255:0] input_199;
    input [255:0] input_200;
    input [255:0] input_201;
    input [255:0] input_202;
    input [255:0] input_203;
    input [255:0] input_204;
    input [255:0] input_205;
    input [255:0] input_206;
    input [255:0] input_207;
    input [255:0] input_208;
    input [255:0] input_209;
    input [255:0] input_210;
    input [255:0] input_211;
    input [255:0] input_212;
    input [255:0] input_213;
    input [255:0] input_214;
    input [255:0] input_215;
    input [255:0] input_216;
    input [255:0] input_217;
    input [255:0] input_218;
    input [255:0] input_219;
    input [255:0] input_220;
    input [255:0] input_221;
    input [255:0] input_222;
    input [255:0] input_223;
    input [255:0] input_224;
    input [255:0] input_225;
    input [255:0] input_226;
    input [255:0] input_227;
    input [255:0] input_228;
    input [255:0] input_229;
    input [255:0] input_230;
    input [255:0] input_231;
    input [255:0] input_232;
    input [255:0] input_233;
    input [255:0] input_234;
    input [255:0] input_235;
    input [255:0] input_236;
    input [255:0] input_237;
    input [255:0] input_238;
    input [255:0] input_239;
    input [255:0] input_240;
    input [255:0] input_241;
    input [255:0] input_242;
    input [255:0] input_243;
    input [255:0] input_244;
    input [255:0] input_245;
    input [255:0] input_246;
    input [255:0] input_247;
    input [255:0] input_248;
    input [255:0] input_249;
    input [255:0] input_250;
    input [255:0] input_251;
    input [255:0] input_252;
    input [255:0] input_253;
    input [255:0] input_254;
    input [255:0] input_255;
    input [7:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      8'b00000000 : begin
        result = input_0;
      end
      8'b00000001 : begin
        result = input_1;
      end
      8'b00000010 : begin
        result = input_2;
      end
      8'b00000011 : begin
        result = input_3;
      end
      8'b00000100 : begin
        result = input_4;
      end
      8'b00000101 : begin
        result = input_5;
      end
      8'b00000110 : begin
        result = input_6;
      end
      8'b00000111 : begin
        result = input_7;
      end
      8'b00001000 : begin
        result = input_8;
      end
      8'b00001001 : begin
        result = input_9;
      end
      8'b00001010 : begin
        result = input_10;
      end
      8'b00001011 : begin
        result = input_11;
      end
      8'b00001100 : begin
        result = input_12;
      end
      8'b00001101 : begin
        result = input_13;
      end
      8'b00001110 : begin
        result = input_14;
      end
      8'b00001111 : begin
        result = input_15;
      end
      8'b00010000 : begin
        result = input_16;
      end
      8'b00010001 : begin
        result = input_17;
      end
      8'b00010010 : begin
        result = input_18;
      end
      8'b00010011 : begin
        result = input_19;
      end
      8'b00010100 : begin
        result = input_20;
      end
      8'b00010101 : begin
        result = input_21;
      end
      8'b00010110 : begin
        result = input_22;
      end
      8'b00010111 : begin
        result = input_23;
      end
      8'b00011000 : begin
        result = input_24;
      end
      8'b00011001 : begin
        result = input_25;
      end
      8'b00011010 : begin
        result = input_26;
      end
      8'b00011011 : begin
        result = input_27;
      end
      8'b00011100 : begin
        result = input_28;
      end
      8'b00011101 : begin
        result = input_29;
      end
      8'b00011110 : begin
        result = input_30;
      end
      8'b00011111 : begin
        result = input_31;
      end
      8'b00100000 : begin
        result = input_32;
      end
      8'b00100001 : begin
        result = input_33;
      end
      8'b00100010 : begin
        result = input_34;
      end
      8'b00100011 : begin
        result = input_35;
      end
      8'b00100100 : begin
        result = input_36;
      end
      8'b00100101 : begin
        result = input_37;
      end
      8'b00100110 : begin
        result = input_38;
      end
      8'b00100111 : begin
        result = input_39;
      end
      8'b00101000 : begin
        result = input_40;
      end
      8'b00101001 : begin
        result = input_41;
      end
      8'b00101010 : begin
        result = input_42;
      end
      8'b00101011 : begin
        result = input_43;
      end
      8'b00101100 : begin
        result = input_44;
      end
      8'b00101101 : begin
        result = input_45;
      end
      8'b00101110 : begin
        result = input_46;
      end
      8'b00101111 : begin
        result = input_47;
      end
      8'b00110000 : begin
        result = input_48;
      end
      8'b00110001 : begin
        result = input_49;
      end
      8'b00110010 : begin
        result = input_50;
      end
      8'b00110011 : begin
        result = input_51;
      end
      8'b00110100 : begin
        result = input_52;
      end
      8'b00110101 : begin
        result = input_53;
      end
      8'b00110110 : begin
        result = input_54;
      end
      8'b00110111 : begin
        result = input_55;
      end
      8'b00111000 : begin
        result = input_56;
      end
      8'b00111001 : begin
        result = input_57;
      end
      8'b00111010 : begin
        result = input_58;
      end
      8'b00111011 : begin
        result = input_59;
      end
      8'b00111100 : begin
        result = input_60;
      end
      8'b00111101 : begin
        result = input_61;
      end
      8'b00111110 : begin
        result = input_62;
      end
      8'b00111111 : begin
        result = input_63;
      end
      8'b01000000 : begin
        result = input_64;
      end
      8'b01000001 : begin
        result = input_65;
      end
      8'b01000010 : begin
        result = input_66;
      end
      8'b01000011 : begin
        result = input_67;
      end
      8'b01000100 : begin
        result = input_68;
      end
      8'b01000101 : begin
        result = input_69;
      end
      8'b01000110 : begin
        result = input_70;
      end
      8'b01000111 : begin
        result = input_71;
      end
      8'b01001000 : begin
        result = input_72;
      end
      8'b01001001 : begin
        result = input_73;
      end
      8'b01001010 : begin
        result = input_74;
      end
      8'b01001011 : begin
        result = input_75;
      end
      8'b01001100 : begin
        result = input_76;
      end
      8'b01001101 : begin
        result = input_77;
      end
      8'b01001110 : begin
        result = input_78;
      end
      8'b01001111 : begin
        result = input_79;
      end
      8'b01010000 : begin
        result = input_80;
      end
      8'b01010001 : begin
        result = input_81;
      end
      8'b01010010 : begin
        result = input_82;
      end
      8'b01010011 : begin
        result = input_83;
      end
      8'b01010100 : begin
        result = input_84;
      end
      8'b01010101 : begin
        result = input_85;
      end
      8'b01010110 : begin
        result = input_86;
      end
      8'b01010111 : begin
        result = input_87;
      end
      8'b01011000 : begin
        result = input_88;
      end
      8'b01011001 : begin
        result = input_89;
      end
      8'b01011010 : begin
        result = input_90;
      end
      8'b01011011 : begin
        result = input_91;
      end
      8'b01011100 : begin
        result = input_92;
      end
      8'b01011101 : begin
        result = input_93;
      end
      8'b01011110 : begin
        result = input_94;
      end
      8'b01011111 : begin
        result = input_95;
      end
      8'b01100000 : begin
        result = input_96;
      end
      8'b01100001 : begin
        result = input_97;
      end
      8'b01100010 : begin
        result = input_98;
      end
      8'b01100011 : begin
        result = input_99;
      end
      8'b01100100 : begin
        result = input_100;
      end
      8'b01100101 : begin
        result = input_101;
      end
      8'b01100110 : begin
        result = input_102;
      end
      8'b01100111 : begin
        result = input_103;
      end
      8'b01101000 : begin
        result = input_104;
      end
      8'b01101001 : begin
        result = input_105;
      end
      8'b01101010 : begin
        result = input_106;
      end
      8'b01101011 : begin
        result = input_107;
      end
      8'b01101100 : begin
        result = input_108;
      end
      8'b01101101 : begin
        result = input_109;
      end
      8'b01101110 : begin
        result = input_110;
      end
      8'b01101111 : begin
        result = input_111;
      end
      8'b01110000 : begin
        result = input_112;
      end
      8'b01110001 : begin
        result = input_113;
      end
      8'b01110010 : begin
        result = input_114;
      end
      8'b01110011 : begin
        result = input_115;
      end
      8'b01110100 : begin
        result = input_116;
      end
      8'b01110101 : begin
        result = input_117;
      end
      8'b01110110 : begin
        result = input_118;
      end
      8'b01110111 : begin
        result = input_119;
      end
      8'b01111000 : begin
        result = input_120;
      end
      8'b01111001 : begin
        result = input_121;
      end
      8'b01111010 : begin
        result = input_122;
      end
      8'b01111011 : begin
        result = input_123;
      end
      8'b01111100 : begin
        result = input_124;
      end
      8'b01111101 : begin
        result = input_125;
      end
      8'b01111110 : begin
        result = input_126;
      end
      8'b01111111 : begin
        result = input_127;
      end
      8'b10000000 : begin
        result = input_128;
      end
      8'b10000001 : begin
        result = input_129;
      end
      8'b10000010 : begin
        result = input_130;
      end
      8'b10000011 : begin
        result = input_131;
      end
      8'b10000100 : begin
        result = input_132;
      end
      8'b10000101 : begin
        result = input_133;
      end
      8'b10000110 : begin
        result = input_134;
      end
      8'b10000111 : begin
        result = input_135;
      end
      8'b10001000 : begin
        result = input_136;
      end
      8'b10001001 : begin
        result = input_137;
      end
      8'b10001010 : begin
        result = input_138;
      end
      8'b10001011 : begin
        result = input_139;
      end
      8'b10001100 : begin
        result = input_140;
      end
      8'b10001101 : begin
        result = input_141;
      end
      8'b10001110 : begin
        result = input_142;
      end
      8'b10001111 : begin
        result = input_143;
      end
      8'b10010000 : begin
        result = input_144;
      end
      8'b10010001 : begin
        result = input_145;
      end
      8'b10010010 : begin
        result = input_146;
      end
      8'b10010011 : begin
        result = input_147;
      end
      8'b10010100 : begin
        result = input_148;
      end
      8'b10010101 : begin
        result = input_149;
      end
      8'b10010110 : begin
        result = input_150;
      end
      8'b10010111 : begin
        result = input_151;
      end
      8'b10011000 : begin
        result = input_152;
      end
      8'b10011001 : begin
        result = input_153;
      end
      8'b10011010 : begin
        result = input_154;
      end
      8'b10011011 : begin
        result = input_155;
      end
      8'b10011100 : begin
        result = input_156;
      end
      8'b10011101 : begin
        result = input_157;
      end
      8'b10011110 : begin
        result = input_158;
      end
      8'b10011111 : begin
        result = input_159;
      end
      8'b10100000 : begin
        result = input_160;
      end
      8'b10100001 : begin
        result = input_161;
      end
      8'b10100010 : begin
        result = input_162;
      end
      8'b10100011 : begin
        result = input_163;
      end
      8'b10100100 : begin
        result = input_164;
      end
      8'b10100101 : begin
        result = input_165;
      end
      8'b10100110 : begin
        result = input_166;
      end
      8'b10100111 : begin
        result = input_167;
      end
      8'b10101000 : begin
        result = input_168;
      end
      8'b10101001 : begin
        result = input_169;
      end
      8'b10101010 : begin
        result = input_170;
      end
      8'b10101011 : begin
        result = input_171;
      end
      8'b10101100 : begin
        result = input_172;
      end
      8'b10101101 : begin
        result = input_173;
      end
      8'b10101110 : begin
        result = input_174;
      end
      8'b10101111 : begin
        result = input_175;
      end
      8'b10110000 : begin
        result = input_176;
      end
      8'b10110001 : begin
        result = input_177;
      end
      8'b10110010 : begin
        result = input_178;
      end
      8'b10110011 : begin
        result = input_179;
      end
      8'b10110100 : begin
        result = input_180;
      end
      8'b10110101 : begin
        result = input_181;
      end
      8'b10110110 : begin
        result = input_182;
      end
      8'b10110111 : begin
        result = input_183;
      end
      8'b10111000 : begin
        result = input_184;
      end
      8'b10111001 : begin
        result = input_185;
      end
      8'b10111010 : begin
        result = input_186;
      end
      8'b10111011 : begin
        result = input_187;
      end
      8'b10111100 : begin
        result = input_188;
      end
      8'b10111101 : begin
        result = input_189;
      end
      8'b10111110 : begin
        result = input_190;
      end
      8'b10111111 : begin
        result = input_191;
      end
      8'b11000000 : begin
        result = input_192;
      end
      8'b11000001 : begin
        result = input_193;
      end
      8'b11000010 : begin
        result = input_194;
      end
      8'b11000011 : begin
        result = input_195;
      end
      8'b11000100 : begin
        result = input_196;
      end
      8'b11000101 : begin
        result = input_197;
      end
      8'b11000110 : begin
        result = input_198;
      end
      8'b11000111 : begin
        result = input_199;
      end
      8'b11001000 : begin
        result = input_200;
      end
      8'b11001001 : begin
        result = input_201;
      end
      8'b11001010 : begin
        result = input_202;
      end
      8'b11001011 : begin
        result = input_203;
      end
      8'b11001100 : begin
        result = input_204;
      end
      8'b11001101 : begin
        result = input_205;
      end
      8'b11001110 : begin
        result = input_206;
      end
      8'b11001111 : begin
        result = input_207;
      end
      8'b11010000 : begin
        result = input_208;
      end
      8'b11010001 : begin
        result = input_209;
      end
      8'b11010010 : begin
        result = input_210;
      end
      8'b11010011 : begin
        result = input_211;
      end
      8'b11010100 : begin
        result = input_212;
      end
      8'b11010101 : begin
        result = input_213;
      end
      8'b11010110 : begin
        result = input_214;
      end
      8'b11010111 : begin
        result = input_215;
      end
      8'b11011000 : begin
        result = input_216;
      end
      8'b11011001 : begin
        result = input_217;
      end
      8'b11011010 : begin
        result = input_218;
      end
      8'b11011011 : begin
        result = input_219;
      end
      8'b11011100 : begin
        result = input_220;
      end
      8'b11011101 : begin
        result = input_221;
      end
      8'b11011110 : begin
        result = input_222;
      end
      8'b11011111 : begin
        result = input_223;
      end
      8'b11100000 : begin
        result = input_224;
      end
      8'b11100001 : begin
        result = input_225;
      end
      8'b11100010 : begin
        result = input_226;
      end
      8'b11100011 : begin
        result = input_227;
      end
      8'b11100100 : begin
        result = input_228;
      end
      8'b11100101 : begin
        result = input_229;
      end
      8'b11100110 : begin
        result = input_230;
      end
      8'b11100111 : begin
        result = input_231;
      end
      8'b11101000 : begin
        result = input_232;
      end
      8'b11101001 : begin
        result = input_233;
      end
      8'b11101010 : begin
        result = input_234;
      end
      8'b11101011 : begin
        result = input_235;
      end
      8'b11101100 : begin
        result = input_236;
      end
      8'b11101101 : begin
        result = input_237;
      end
      8'b11101110 : begin
        result = input_238;
      end
      8'b11101111 : begin
        result = input_239;
      end
      8'b11110000 : begin
        result = input_240;
      end
      8'b11110001 : begin
        result = input_241;
      end
      8'b11110010 : begin
        result = input_242;
      end
      8'b11110011 : begin
        result = input_243;
      end
      8'b11110100 : begin
        result = input_244;
      end
      8'b11110101 : begin
        result = input_245;
      end
      8'b11110110 : begin
        result = input_246;
      end
      8'b11110111 : begin
        result = input_247;
      end
      8'b11111000 : begin
        result = input_248;
      end
      8'b11111001 : begin
        result = input_249;
      end
      8'b11111010 : begin
        result = input_250;
      end
      8'b11111011 : begin
        result = input_251;
      end
      8'b11111100 : begin
        result = input_252;
      end
      8'b11111101 : begin
        result = input_253;
      end
      8'b11111110 : begin
        result = input_254;
      end
      default : begin
        result = input_255;
      end
    endcase
    MUX_v_256_256_2 = result;
  end
  endfunction


  function automatic [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input  sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [35:0] MUX_v_36_2_2;
    input [35:0] input_0;
    input [35:0] input_1;
    input  sel;
    reg [35:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_36_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [10:0] signext_11_1;
    input  vector;
  begin
    signext_11_1= {{10{vector}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input  vector;
  begin
    signext_4_1= {{3{vector}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input  vector;
  begin
    signext_7_1= {{6{vector}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [35:0] conv_u2s_35_36 ;
    input [34:0]  vector ;
  begin
    conv_u2s_35_36 =  {1'b0, vector};
  end
  endfunction


  function automatic [34:0] conv_u2u_34_35 ;
    input [33:0]  vector ;
  begin
    conv_u2u_34_35 = {1'b0, vector};
  end
  endfunction


  function automatic [35:0] conv_u2u_34_36 ;
    input [33:0]  vector ;
  begin
    conv_u2u_34_36 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore
// ------------------------------------------------------------------


module PECore (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [265:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [312:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [255:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  wire [255:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  wire [255:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  wire [255:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  wire [255:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  wire [255:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  wire [255:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  wire [255:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  wire [255:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  wire [255:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  wire [255:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  wire [255:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  wire [255:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  wire [255:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  wire [255:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  wire [255:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  wire [255:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_c;
  wire Datapath_for_4_ProductSum_for_acc_9_cmp_en;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_b;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_c;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_d;
  wire Datapath_for_4_ProductSum_for_acc_9_cmp_1_en;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_1_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_b;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_c;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_d;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_2_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_b;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_c;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_d;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_3_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_b;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_c;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_d;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_4_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_b;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_c;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_d;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_5_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_b;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_c;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_d;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_6_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_b;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_c;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_d;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_7_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_16_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_17_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_18_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_19_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_20_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_21_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_22_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_23_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_24_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_25_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_26_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_27_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_28_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_29_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_30_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_31_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_32_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_33_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_34_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_35_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_36_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_37_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_38_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_39_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_40_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_41_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_42_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_43_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_44_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_45_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_46_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_47_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_48_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_49_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_50_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_51_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_52_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_53_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_54_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_55_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_56_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_57_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_58_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_59_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_60_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_61_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_62_z;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_a;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_c;
  wire [33:0] Datapath_for_4_ProductSum_for_acc_9_cmp_63_z;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_clken;
  wire [255:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_we;
  wire [255:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_clken;
  wire [255:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_we;
  wire [255:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_clken;
  wire [255:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_we;
  wire [255:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_clken;
  wire [255:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_we;
  wire [255:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_clken;
  wire [255:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_we;
  wire [255:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_clken;
  wire [255:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_we;
  wire [255:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_clken;
  wire [255:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_we;
  wire [255:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_clken;
  wire [255:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_we;
  wire [255:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_iff;
  wire [15:0] Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_1 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_1_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_1_b),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_1_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_1_d),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_1_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_2 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_2_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_2_b),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_2_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_2_d),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_2_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_3 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_3_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_3_b),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_3_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_3_d),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_3_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_4 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_4_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_4_b),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_4_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_4_d),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_4_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_5 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_5_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_5_b),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_5_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_5_d),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_5_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_6 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_6_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_6_b),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_6_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_6_d),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_6_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_7 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_7_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_7_b),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_7_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_7_d),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_7_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_8 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_8_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_8_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_8_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_9 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_9_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_9_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_9_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_10 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_10_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_10_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_10_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_11 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_11_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_11_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_11_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_12 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_12_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_12_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_12_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_13 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_13_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_13_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_13_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_14 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_14_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_14_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_14_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_15 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_15_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_15_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_15_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_16 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_16_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_16_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_16_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_17 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_17_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_17_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_17_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_18 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_18_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_18_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_18_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_19 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_19_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_19_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_19_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_20 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_20_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_20_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_20_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_21 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_21_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_21_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_21_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_22 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_22_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_22_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_22_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_23 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_23_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_23_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_23_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_24 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_24_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_24_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_24_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_25 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_25_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_25_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_25_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_26 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_26_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_26_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_26_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_27 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_27_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_27_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_27_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_28 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_28_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_28_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_28_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_29 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_29_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_29_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_29_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_30 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_30_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_30_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_30_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_31 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_31_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_31_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_31_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_32 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_32_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_32_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_32_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_33 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_33_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_33_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_33_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_34 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_34_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_34_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_34_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_35 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_35_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_35_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_35_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_36 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_36_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_36_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_36_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_37 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_37_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_37_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_37_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_38 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_38_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_38_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_38_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_39 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_39_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_39_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_39_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_40 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_40_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_40_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_40_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_41 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_41_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_41_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_41_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_42 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_42_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_42_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_42_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_43 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_43_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_43_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_43_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_44 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_44_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_44_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_44_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_45 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_45_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_45_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_45_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_46 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_46_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_46_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_46_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_47 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_47_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_47_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_47_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_48 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_48_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_48_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_48_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_49 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_49_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_49_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_49_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_50 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_50_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_50_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_50_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_51 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_51_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_51_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_51_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_52 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_52_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_52_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_52_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_53 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_53_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_53_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_53_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_54 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_54_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_54_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_54_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_55 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_55_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_55_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_55_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_56 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_56_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_56_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_56_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_57 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_57_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_57_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_57_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_58 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_58_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_58_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_58_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_59 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_59_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_59_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_59_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_60 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_60_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_60_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_60_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_61 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_61_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_61_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_61_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_62 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_62_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_62_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_62_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd16),
  .signd_a(32'sd0),
  .width_b(32'sd16),
  .signd_b(32'sd0),
  .width_c(32'sd16),
  .signd_c(32'sd0),
  .width_d(32'sd16),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd34),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_9_cmp_63 (
      .a(Datapath_for_4_ProductSum_for_acc_9_cmp_63_a),
      .b(Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_9_cmp_63_c),
      .d(Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_9_cmp_63_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd256),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd256),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd256),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd256),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd256),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd256),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd256),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd256),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_256_4096_1_4096_256_1_gen
      weight_mem_banks_bank_a0_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_256_4096_1_4096_256_1_gen
      weight_mem_banks_bank_a0_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_256_4096_1_4096_256_1_gen
      weight_mem_banks_bank_a0_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_256_4096_1_4096_256_1_gen
      weight_mem_banks_bank_a0_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_256_4096_1_4096_256_1_gen
      weight_mem_banks_bank_a1_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_256_4096_1_4096_256_1_gen
      weight_mem_banks_bank_a1_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_256_4096_1_4096_256_1_gen
      weight_mem_banks_bank_a1_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_256_4096_1_4096_256_1_gen
      weight_mem_banks_bank_a1_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_PECoreRun PECore_PECoreRun_inst (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_a(Datapath_for_4_ProductSum_for_acc_9_cmp_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_c(Datapath_for_4_ProductSum_for_acc_9_cmp_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_en(Datapath_for_4_ProductSum_for_acc_9_cmp_en),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_z(Datapath_for_4_ProductSum_for_acc_9_cmp_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_a(Datapath_for_4_ProductSum_for_acc_9_cmp_1_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_b(Datapath_for_4_ProductSum_for_acc_9_cmp_1_b),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_c(Datapath_for_4_ProductSum_for_acc_9_cmp_1_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_d(Datapath_for_4_ProductSum_for_acc_9_cmp_1_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_en(Datapath_for_4_ProductSum_for_acc_9_cmp_1_en),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_1_z(Datapath_for_4_ProductSum_for_acc_9_cmp_1_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_a(Datapath_for_4_ProductSum_for_acc_9_cmp_2_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_b(Datapath_for_4_ProductSum_for_acc_9_cmp_2_b),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_c(Datapath_for_4_ProductSum_for_acc_9_cmp_2_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_d(Datapath_for_4_ProductSum_for_acc_9_cmp_2_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_2_z(Datapath_for_4_ProductSum_for_acc_9_cmp_2_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_a(Datapath_for_4_ProductSum_for_acc_9_cmp_3_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_b(Datapath_for_4_ProductSum_for_acc_9_cmp_3_b),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_c(Datapath_for_4_ProductSum_for_acc_9_cmp_3_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_d(Datapath_for_4_ProductSum_for_acc_9_cmp_3_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_3_z(Datapath_for_4_ProductSum_for_acc_9_cmp_3_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_a(Datapath_for_4_ProductSum_for_acc_9_cmp_4_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_b(Datapath_for_4_ProductSum_for_acc_9_cmp_4_b),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_c(Datapath_for_4_ProductSum_for_acc_9_cmp_4_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_d(Datapath_for_4_ProductSum_for_acc_9_cmp_4_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_4_z(Datapath_for_4_ProductSum_for_acc_9_cmp_4_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_a(Datapath_for_4_ProductSum_for_acc_9_cmp_5_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_b(Datapath_for_4_ProductSum_for_acc_9_cmp_5_b),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_c(Datapath_for_4_ProductSum_for_acc_9_cmp_5_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_d(Datapath_for_4_ProductSum_for_acc_9_cmp_5_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_5_z(Datapath_for_4_ProductSum_for_acc_9_cmp_5_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_a(Datapath_for_4_ProductSum_for_acc_9_cmp_6_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_b(Datapath_for_4_ProductSum_for_acc_9_cmp_6_b),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_c(Datapath_for_4_ProductSum_for_acc_9_cmp_6_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_d(Datapath_for_4_ProductSum_for_acc_9_cmp_6_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_6_z(Datapath_for_4_ProductSum_for_acc_9_cmp_6_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_a(Datapath_for_4_ProductSum_for_acc_9_cmp_7_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_b(Datapath_for_4_ProductSum_for_acc_9_cmp_7_b),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_c(Datapath_for_4_ProductSum_for_acc_9_cmp_7_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_d(Datapath_for_4_ProductSum_for_acc_9_cmp_7_d),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_7_z(Datapath_for_4_ProductSum_for_acc_9_cmp_7_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_a(Datapath_for_4_ProductSum_for_acc_9_cmp_8_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_c(Datapath_for_4_ProductSum_for_acc_9_cmp_8_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_z(Datapath_for_4_ProductSum_for_acc_9_cmp_8_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_9_a(Datapath_for_4_ProductSum_for_acc_9_cmp_9_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_9_c(Datapath_for_4_ProductSum_for_acc_9_cmp_9_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_9_z(Datapath_for_4_ProductSum_for_acc_9_cmp_9_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_10_a(Datapath_for_4_ProductSum_for_acc_9_cmp_10_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_10_c(Datapath_for_4_ProductSum_for_acc_9_cmp_10_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_10_z(Datapath_for_4_ProductSum_for_acc_9_cmp_10_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_11_a(Datapath_for_4_ProductSum_for_acc_9_cmp_11_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_11_c(Datapath_for_4_ProductSum_for_acc_9_cmp_11_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_11_z(Datapath_for_4_ProductSum_for_acc_9_cmp_11_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_12_a(Datapath_for_4_ProductSum_for_acc_9_cmp_12_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_12_c(Datapath_for_4_ProductSum_for_acc_9_cmp_12_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_12_z(Datapath_for_4_ProductSum_for_acc_9_cmp_12_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_13_a(Datapath_for_4_ProductSum_for_acc_9_cmp_13_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_13_c(Datapath_for_4_ProductSum_for_acc_9_cmp_13_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_13_z(Datapath_for_4_ProductSum_for_acc_9_cmp_13_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_14_a(Datapath_for_4_ProductSum_for_acc_9_cmp_14_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_14_c(Datapath_for_4_ProductSum_for_acc_9_cmp_14_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_14_z(Datapath_for_4_ProductSum_for_acc_9_cmp_14_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_15_a(Datapath_for_4_ProductSum_for_acc_9_cmp_15_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_15_c(Datapath_for_4_ProductSum_for_acc_9_cmp_15_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_15_z(Datapath_for_4_ProductSum_for_acc_9_cmp_15_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_16_a(Datapath_for_4_ProductSum_for_acc_9_cmp_16_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_16_c(Datapath_for_4_ProductSum_for_acc_9_cmp_16_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_16_z(Datapath_for_4_ProductSum_for_acc_9_cmp_16_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_17_a(Datapath_for_4_ProductSum_for_acc_9_cmp_17_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_17_c(Datapath_for_4_ProductSum_for_acc_9_cmp_17_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_17_z(Datapath_for_4_ProductSum_for_acc_9_cmp_17_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_18_a(Datapath_for_4_ProductSum_for_acc_9_cmp_18_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_18_c(Datapath_for_4_ProductSum_for_acc_9_cmp_18_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_18_z(Datapath_for_4_ProductSum_for_acc_9_cmp_18_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_19_a(Datapath_for_4_ProductSum_for_acc_9_cmp_19_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_19_c(Datapath_for_4_ProductSum_for_acc_9_cmp_19_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_19_z(Datapath_for_4_ProductSum_for_acc_9_cmp_19_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_20_a(Datapath_for_4_ProductSum_for_acc_9_cmp_20_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_20_c(Datapath_for_4_ProductSum_for_acc_9_cmp_20_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_20_z(Datapath_for_4_ProductSum_for_acc_9_cmp_20_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_21_a(Datapath_for_4_ProductSum_for_acc_9_cmp_21_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_21_c(Datapath_for_4_ProductSum_for_acc_9_cmp_21_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_21_z(Datapath_for_4_ProductSum_for_acc_9_cmp_21_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_22_a(Datapath_for_4_ProductSum_for_acc_9_cmp_22_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_22_c(Datapath_for_4_ProductSum_for_acc_9_cmp_22_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_22_z(Datapath_for_4_ProductSum_for_acc_9_cmp_22_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_23_a(Datapath_for_4_ProductSum_for_acc_9_cmp_23_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_23_c(Datapath_for_4_ProductSum_for_acc_9_cmp_23_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_23_z(Datapath_for_4_ProductSum_for_acc_9_cmp_23_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_24_a(Datapath_for_4_ProductSum_for_acc_9_cmp_24_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_24_c(Datapath_for_4_ProductSum_for_acc_9_cmp_24_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_24_z(Datapath_for_4_ProductSum_for_acc_9_cmp_24_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_25_a(Datapath_for_4_ProductSum_for_acc_9_cmp_25_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_25_c(Datapath_for_4_ProductSum_for_acc_9_cmp_25_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_25_z(Datapath_for_4_ProductSum_for_acc_9_cmp_25_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_26_a(Datapath_for_4_ProductSum_for_acc_9_cmp_26_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_26_c(Datapath_for_4_ProductSum_for_acc_9_cmp_26_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_26_z(Datapath_for_4_ProductSum_for_acc_9_cmp_26_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_27_a(Datapath_for_4_ProductSum_for_acc_9_cmp_27_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_27_c(Datapath_for_4_ProductSum_for_acc_9_cmp_27_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_27_z(Datapath_for_4_ProductSum_for_acc_9_cmp_27_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_28_a(Datapath_for_4_ProductSum_for_acc_9_cmp_28_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_28_c(Datapath_for_4_ProductSum_for_acc_9_cmp_28_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_28_z(Datapath_for_4_ProductSum_for_acc_9_cmp_28_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_29_a(Datapath_for_4_ProductSum_for_acc_9_cmp_29_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_29_c(Datapath_for_4_ProductSum_for_acc_9_cmp_29_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_29_z(Datapath_for_4_ProductSum_for_acc_9_cmp_29_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_30_a(Datapath_for_4_ProductSum_for_acc_9_cmp_30_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_30_c(Datapath_for_4_ProductSum_for_acc_9_cmp_30_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_30_z(Datapath_for_4_ProductSum_for_acc_9_cmp_30_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_31_a(Datapath_for_4_ProductSum_for_acc_9_cmp_31_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_31_c(Datapath_for_4_ProductSum_for_acc_9_cmp_31_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_31_z(Datapath_for_4_ProductSum_for_acc_9_cmp_31_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_32_a(Datapath_for_4_ProductSum_for_acc_9_cmp_32_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_32_c(Datapath_for_4_ProductSum_for_acc_9_cmp_32_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_32_z(Datapath_for_4_ProductSum_for_acc_9_cmp_32_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_33_a(Datapath_for_4_ProductSum_for_acc_9_cmp_33_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_33_c(Datapath_for_4_ProductSum_for_acc_9_cmp_33_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_33_z(Datapath_for_4_ProductSum_for_acc_9_cmp_33_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_34_a(Datapath_for_4_ProductSum_for_acc_9_cmp_34_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_34_c(Datapath_for_4_ProductSum_for_acc_9_cmp_34_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_34_z(Datapath_for_4_ProductSum_for_acc_9_cmp_34_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_35_a(Datapath_for_4_ProductSum_for_acc_9_cmp_35_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_35_c(Datapath_for_4_ProductSum_for_acc_9_cmp_35_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_35_z(Datapath_for_4_ProductSum_for_acc_9_cmp_35_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_36_a(Datapath_for_4_ProductSum_for_acc_9_cmp_36_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_36_c(Datapath_for_4_ProductSum_for_acc_9_cmp_36_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_36_z(Datapath_for_4_ProductSum_for_acc_9_cmp_36_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_37_a(Datapath_for_4_ProductSum_for_acc_9_cmp_37_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_37_c(Datapath_for_4_ProductSum_for_acc_9_cmp_37_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_37_z(Datapath_for_4_ProductSum_for_acc_9_cmp_37_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_38_a(Datapath_for_4_ProductSum_for_acc_9_cmp_38_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_38_c(Datapath_for_4_ProductSum_for_acc_9_cmp_38_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_38_z(Datapath_for_4_ProductSum_for_acc_9_cmp_38_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_39_a(Datapath_for_4_ProductSum_for_acc_9_cmp_39_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_39_c(Datapath_for_4_ProductSum_for_acc_9_cmp_39_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_39_z(Datapath_for_4_ProductSum_for_acc_9_cmp_39_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_40_a(Datapath_for_4_ProductSum_for_acc_9_cmp_40_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_40_c(Datapath_for_4_ProductSum_for_acc_9_cmp_40_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_40_z(Datapath_for_4_ProductSum_for_acc_9_cmp_40_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_41_a(Datapath_for_4_ProductSum_for_acc_9_cmp_41_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_41_c(Datapath_for_4_ProductSum_for_acc_9_cmp_41_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_41_z(Datapath_for_4_ProductSum_for_acc_9_cmp_41_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_42_a(Datapath_for_4_ProductSum_for_acc_9_cmp_42_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_42_c(Datapath_for_4_ProductSum_for_acc_9_cmp_42_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_42_z(Datapath_for_4_ProductSum_for_acc_9_cmp_42_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_43_a(Datapath_for_4_ProductSum_for_acc_9_cmp_43_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_43_c(Datapath_for_4_ProductSum_for_acc_9_cmp_43_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_43_z(Datapath_for_4_ProductSum_for_acc_9_cmp_43_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_44_a(Datapath_for_4_ProductSum_for_acc_9_cmp_44_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_44_c(Datapath_for_4_ProductSum_for_acc_9_cmp_44_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_44_z(Datapath_for_4_ProductSum_for_acc_9_cmp_44_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_45_a(Datapath_for_4_ProductSum_for_acc_9_cmp_45_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_45_c(Datapath_for_4_ProductSum_for_acc_9_cmp_45_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_45_z(Datapath_for_4_ProductSum_for_acc_9_cmp_45_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_46_a(Datapath_for_4_ProductSum_for_acc_9_cmp_46_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_46_c(Datapath_for_4_ProductSum_for_acc_9_cmp_46_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_46_z(Datapath_for_4_ProductSum_for_acc_9_cmp_46_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_47_a(Datapath_for_4_ProductSum_for_acc_9_cmp_47_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_47_c(Datapath_for_4_ProductSum_for_acc_9_cmp_47_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_47_z(Datapath_for_4_ProductSum_for_acc_9_cmp_47_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_48_a(Datapath_for_4_ProductSum_for_acc_9_cmp_48_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_48_c(Datapath_for_4_ProductSum_for_acc_9_cmp_48_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_48_z(Datapath_for_4_ProductSum_for_acc_9_cmp_48_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_49_a(Datapath_for_4_ProductSum_for_acc_9_cmp_49_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_49_c(Datapath_for_4_ProductSum_for_acc_9_cmp_49_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_49_z(Datapath_for_4_ProductSum_for_acc_9_cmp_49_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_50_a(Datapath_for_4_ProductSum_for_acc_9_cmp_50_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_50_c(Datapath_for_4_ProductSum_for_acc_9_cmp_50_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_50_z(Datapath_for_4_ProductSum_for_acc_9_cmp_50_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_51_a(Datapath_for_4_ProductSum_for_acc_9_cmp_51_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_51_c(Datapath_for_4_ProductSum_for_acc_9_cmp_51_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_51_z(Datapath_for_4_ProductSum_for_acc_9_cmp_51_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_52_a(Datapath_for_4_ProductSum_for_acc_9_cmp_52_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_52_c(Datapath_for_4_ProductSum_for_acc_9_cmp_52_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_52_z(Datapath_for_4_ProductSum_for_acc_9_cmp_52_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_53_a(Datapath_for_4_ProductSum_for_acc_9_cmp_53_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_53_c(Datapath_for_4_ProductSum_for_acc_9_cmp_53_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_53_z(Datapath_for_4_ProductSum_for_acc_9_cmp_53_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_54_a(Datapath_for_4_ProductSum_for_acc_9_cmp_54_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_54_c(Datapath_for_4_ProductSum_for_acc_9_cmp_54_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_54_z(Datapath_for_4_ProductSum_for_acc_9_cmp_54_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_55_a(Datapath_for_4_ProductSum_for_acc_9_cmp_55_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_55_c(Datapath_for_4_ProductSum_for_acc_9_cmp_55_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_55_z(Datapath_for_4_ProductSum_for_acc_9_cmp_55_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_56_a(Datapath_for_4_ProductSum_for_acc_9_cmp_56_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_56_c(Datapath_for_4_ProductSum_for_acc_9_cmp_56_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_56_z(Datapath_for_4_ProductSum_for_acc_9_cmp_56_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_57_a(Datapath_for_4_ProductSum_for_acc_9_cmp_57_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_57_c(Datapath_for_4_ProductSum_for_acc_9_cmp_57_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_57_z(Datapath_for_4_ProductSum_for_acc_9_cmp_57_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_58_a(Datapath_for_4_ProductSum_for_acc_9_cmp_58_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_58_c(Datapath_for_4_ProductSum_for_acc_9_cmp_58_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_58_z(Datapath_for_4_ProductSum_for_acc_9_cmp_58_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_59_a(Datapath_for_4_ProductSum_for_acc_9_cmp_59_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_59_c(Datapath_for_4_ProductSum_for_acc_9_cmp_59_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_59_z(Datapath_for_4_ProductSum_for_acc_9_cmp_59_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_60_a(Datapath_for_4_ProductSum_for_acc_9_cmp_60_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_60_c(Datapath_for_4_ProductSum_for_acc_9_cmp_60_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_60_z(Datapath_for_4_ProductSum_for_acc_9_cmp_60_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_61_a(Datapath_for_4_ProductSum_for_acc_9_cmp_61_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_61_c(Datapath_for_4_ProductSum_for_acc_9_cmp_61_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_61_z(Datapath_for_4_ProductSum_for_acc_9_cmp_61_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_62_a(Datapath_for_4_ProductSum_for_acc_9_cmp_62_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_62_c(Datapath_for_4_ProductSum_for_acc_9_cmp_62_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_62_z(Datapath_for_4_ProductSum_for_acc_9_cmp_62_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_63_a(Datapath_for_4_ProductSum_for_acc_9_cmp_63_a),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_63_c(Datapath_for_4_ProductSum_for_acc_9_cmp_63_c),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_63_z(Datapath_for_4_ProductSum_for_acc_9_cmp_63_z),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_8_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_8_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_9_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_9_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_10_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_10_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_11_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_11_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_12_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_12_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_13_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_13_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_14_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_14_d_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_15_b_iff),
      .Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_pff(Datapath_for_4_ProductSum_for_acc_9_cmp_15_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff)
    );
endmodule



