
//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 01:33:07 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [96:0] this_dat;
  output [63:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [63:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_dat[63:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_dat[87:64];
  wire  nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_dat[96];
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd64)) data_data_rsci (
      .d(nl_data_data_rsci_d[63:0]),
      .z(data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d),
      .z(data_rw_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd154),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [96:0] this_dat;
  output [63:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 01:32:57 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [73:0] this_dat;
  output [63:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [63:0] nl_data_data_data_rsci_d;
  assign nl_data_data_data_rsci_d = this_dat[63:0];
  wire [7:0] nl_data_logical_addr_rsci_d;
  assign nl_data_logical_addr_rsci_d = this_dat[73:66];
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd7),
  .width(32'sd64)) data_data_data_rsci (
      .d(nl_data_data_data_rsci_d[63:0]),
      .z(data_data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd9),
  .width(32'sd8)) data_logical_addr_rsci (
      .d(nl_data_logical_addr_rsci_d[7:0]),
      .z(data_logical_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd11),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd153),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [73:0] this_dat;
  output [63:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_data_rsc_z(data_data_data_rsc_z),
      .data_logical_addr_rsc_z(data_logical_addr_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 01:32:53 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [255:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [15:0] m_data_buf_239_0_lpi_1_dfm_239_224;
  reg [15:0] m_data_buf_239_0_lpi_1_dfm_207_192;
  reg [15:0] m_data_buf_239_0_lpi_1_dfm_175_160;
  reg [15:0] m_data_buf_239_0_lpi_1_dfm_143_128;
  reg [15:0] m_data_buf_239_0_lpi_1_dfm_111_96;
  reg [15:0] m_data_buf_239_0_lpi_1_dfm_79_64;
  reg [15:0] m_data_buf_239_0_lpi_1_dfm_47_32;
  reg [15:0] m_data_buf_239_0_lpi_1_dfm_15_0;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd13),
  .width(32'sd256)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd152),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd156)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = {16'b0000000000000000 , m_data_buf_239_0_lpi_1_dfm_239_224 ,
      16'b0000000000000000 , m_data_buf_239_0_lpi_1_dfm_207_192 , 16'b0000000000000000
      , m_data_buf_239_0_lpi_1_dfm_175_160 , 16'b0000000000000000 , m_data_buf_239_0_lpi_1_dfm_143_128
      , 16'b0000000000000000 , m_data_buf_239_0_lpi_1_dfm_111_96 , 16'b0000000000000000
      , m_data_buf_239_0_lpi_1_dfm_79_64 , 16'b0000000000000000 , m_data_buf_239_0_lpi_1_dfm_47_32
      , 16'b0000000000000000 , m_data_buf_239_0_lpi_1_dfm_15_0};
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_239_0_lpi_1_dfm_239_224 <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_239_0_lpi_1_dfm_239_224 <= m_data_rsci_idat[239:224];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_239_0_lpi_1_dfm_207_192 <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_239_0_lpi_1_dfm_207_192 <= m_data_rsci_idat[207:192];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_239_0_lpi_1_dfm_175_160 <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_239_0_lpi_1_dfm_175_160 <= m_data_rsci_idat[175:160];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_239_0_lpi_1_dfm_143_128 <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_239_0_lpi_1_dfm_143_128 <= m_data_rsci_idat[143:128];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_239_0_lpi_1_dfm_111_96 <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_239_0_lpi_1_dfm_111_96 <= m_data_rsci_idat[111:96];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_239_0_lpi_1_dfm_79_64 <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_239_0_lpi_1_dfm_79_64 <= m_data_rsci_idat[79:64];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_239_0_lpi_1_dfm_47_32 <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_239_0_lpi_1_dfm_47_32 <= m_data_rsci_idat[47:32];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_buf_239_0_lpi_1_dfm_15_0 <= 16'b0000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_buf_239_0_lpi_1_dfm_15_0 <= m_data_rsci_idat[15:0];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 01:32:50 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd15),
  .width(32'sd1)) data_rsci (
      .d(this_dat),
      .z(data_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd17),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd151),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 01:33:03 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [63:0] this_dat;
  reg [63:0] this_dat;
  input [63:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [63:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd18),
  .width(32'sd64)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd150),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd155)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [63:0] this_dat;
  input [63:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_mgc_muladd1_beh.v 
//muladd1
module PECore_mgc_muladd1(a,b,c,cst,d,z);
  // operation is z = a * (b + d) + c + cst
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_cst = 0;
  parameter signd_cst = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_axb = 1;
  parameter add_c = 1;
  parameter add_d = 1;
  parameter use_const = 1;

  function integer is_square_op;
    input integer alen;
  begin
    if (alen > 1) is_square_op = 0;
    else       is_square_op = 1;
  end endfunction

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_cst-1:0] cst; // spyglass disable SYNTH_5121,W240
  input  [width_d-1:0] d;
  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa;
  reg [width_b-signd_b:0] bb;
  reg [width_c-signd_c:0] cc;
  reg [width_d-signd_d:0] dd;
  reg [width_cst-signd_cst:0] cstin;

  localparam width_bd = (width_d) ? 1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b
                                                                          : width_d - signd_d)
                                  : width_b - signd_b;
  localparam is_square = is_square_op(width_a);
  localparam axb_len = (is_square)?width_bd+1+width_bd+1:width_a-signd_a+1+width_bd+1;

  reg [width_bd:0] bd;
  reg [axb_len-1:0] axb;



  // make all inputs signed
  always @(*) aa = signd_a ? a : {1'b0, a};
  always @(*) bb = signd_b ? b : {1'b0, b};
  generate if (width_c != 0) begin
    always @(*) cc = signd_c ? c : {1'b0, c};
  end endgenerate

  generate if (width_d) begin
    if ( !is_square) begin
      (* keep ="true" *) reg [width_d-signd_d:0] d_keep;
      always @(*) d_keep = signd_d ? d : {1'b0, d};
      always @(*) dd = d_keep;
    end else begin
      always @(*) dd = signd_d ? d : {1'b0, d};
    end
  end endgenerate

  always @(*) cstin = signd_cst ? cst : {1'b0, cst};

  // perform pre-adder
  generate
    if (width_d != 0) begin
      if (add_d) begin always @(*)  bd = $signed(bb) + $signed(dd); end
      else       begin always @(*)  bd = $signed(bb) - $signed(dd); end
    end else     begin always @(*)  bd = $signed(bb); end
  endgenerate

  generate
    if (is_square)
      always @(*) axb = $signed(bd) * $signed(bd);
    else
      always @(*) axb = $signed(aa) * $signed(bd);
  endgenerate

  // perform muladd1
  wire [width_z-1:0]  zz;

  generate
    if (use_const) begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc) + $signed(cstin); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc) + $signed(cstin); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb) + $signed(cstin); end else
      if (!add_axb && !add_c && width_c) begin assign zz = $signed(cstin) - $signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb) + $signed(cstin); end else
                                         begin assign zz = $signed(cstin) - $signed(axb); end
    end  else begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb); end else
      if (!add_axb && !add_c && width_c) begin assign zz = -$signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb); end else
                                         begin assign zz = -$signed(axb); end
    end
  endgenerate

  // adjust output
  assign z = zz;
endmodule // mgc_muladd1

//------> ./PECore_mgc_shift_l_beh_v5.v 
module PECore_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./PECore_mgc_mul2add1_pipe_beh.v 
//muladd1
module PECore_mgc_mul2add1_pipe(a,b,b2,c,d,d2,cst,clk,en,a_rst,s_rst,z);
  parameter gentype = 0;
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_b2 = 0;
  parameter signd_b2 = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_d2 = 0;
  parameter signd_d2 = 0;
  parameter width_e = 0;
  parameter signd_e = 0;
  parameter width_z = 0;
  parameter isadd = 1;
  parameter add_b2 = 1;
  parameter add_d2 = 1;
  parameter use_const = 1;
  parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
  parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
  parameter    a_rst_active =  1'b1;  // unused
  parameter    s_rst_active =  1'b1;  // unused
  parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
  parameter integer n_inreg = 32'd0;  // number of input registers

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_b2-1:0] b2; // spyglass disable SYNTH_5121,W240
  input  [width_c-1:0] c;
  input  [width_d-1:0] d;
  input  [width_d2-1:0] d2; // spyglass disable SYNTH_5121,W240
  input  [width_e-1:0] cst; // spyglass disable SYNTH_5121,W240

  input                clk;    // clock
  input                en;     // enable
  input                a_rst;  // spyglass disable SYNTH_5121,W240
  input                s_rst;  // spyglass disable SYNTH_5121,W240

  output [width_z-1:0] z;

  function integer MIN;
    input integer a, b;
  begin
    if (a > b) MIN = b;
    else       MIN = a;
  end endfunction

  function integer f_axb_stages;
    input integer gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d;
  begin
    if (gentype%2==0) begin
      if ((n_inreg > 1) && (width_a>18 | width_b>=19+signd_b | width_c>18 | width_d>=19+signd_d ))
        f_axb_stages = 1;
      else
        f_axb_stages = 0;
    end else begin
      if (n_inreg>1)
        f_axb_stages = 1;
      else
        f_axb_stages = 0;
    end
  end endfunction

  function integer f_cxd_stages;
    input integer gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d;
  begin
    if (gentype%2==0) begin
      f_cxd_stages = 0;
    end else begin
      if (n_inreg>1)
        f_cxd_stages = MIN(n_inreg-1,3);
      else
        f_cxd_stages = 0;
    end
  end endfunction

  function integer f_preadd_stages;
    input integer gentype,n_inreg,width_preaddin;
  begin
    if (gentype%2==0) begin
      f_preadd_stages = 0;
    end else begin
      if (n_inreg>1) begin
        if (width_preaddin>0)
          f_preadd_stages = 1;
        else
          f_preadd_stages = 0;
      end else
        f_preadd_stages = 0;
    end
  end endfunction

  function integer MAX;
    input integer LEFT, RIGHT;
  begin
    if (LEFT > RIGHT) MAX = LEFT;
    else              MAX = RIGHT;
  end endfunction

  function integer PREADDLEN;
    input integer b_len, d_len, width_d;
  begin
    if(width_d>0) PREADDLEN = MAX(b_len,d_len) + 1;
    else        PREADDLEN = b_len;
  end endfunction
  function integer PREADDMULLEN;
    input integer a_len, b_len, d_len, width_d;
  begin
    PREADDMULLEN = a_len + PREADDLEN(b_len,d_len,width_d);
  end endfunction

  localparam axb_stages = f_axb_stages(gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d);
  localparam cxd_stages = f_cxd_stages(gentype,n_inreg,width_a, signd_a,width_b,signd_b,width_c, signd_c,width_d,signd_d);
  localparam preadd_ab_stages = f_preadd_stages(gentype, n_inreg - axb_stages,width_b2);
  localparam preadd_cd_stages = f_preadd_stages(gentype, n_inreg - cxd_stages,width_d2);
  localparam e_stages  = (use_const>1)?n_inreg:0;
  localparam a_stages  = n_inreg - axb_stages;
  localparam b_stages  = n_inreg - axb_stages - preadd_ab_stages;
  localparam c_stages  = n_inreg - cxd_stages;
  localparam d_stages  = n_inreg - cxd_stages - preadd_cd_stages;
  localparam b2_stages  = (width_b2>0)?b_stages:0;
  localparam d2_stages  = (width_d2>0)?d_stages:0;

  localparam a_len    = width_a-signd_a+1;
  localparam b_len    = width_b-signd_b+1;
  localparam b2_len   = width_b2-signd_b2+1;
  localparam c_len    = width_c-signd_c+1;
  localparam d_len    = width_d-signd_d+1;
  localparam d2_len   = width_d2-signd_d2+1;
  localparam e_len    = width_e-signd_e+1;
  localparam bb2_len  = PREADDLEN(b_len, b2_len, width_b2);
  localparam dd2_len  = PREADDLEN(d_len, d2_len, width_d2);
  localparam axb_len  = PREADDMULLEN(a_len, b_len, b2_len, width_b2);
  localparam cxd_len  = PREADDMULLEN(c_len, d_len, d2_len, width_d2);
  localparam z_len    = width_z;

  reg [a_len-1:0]  aa  [a_stages:0];
  reg [b_len-1:0]  bb  [b_stages:0];
  reg [b2_len-1:0] bb2 [b2_stages:0];
  reg [c_len-1:0]  cc  [c_stages:0];
  reg [d_len-1:0]  dd  [d_stages:0];
  reg [d2_len-1:0] dd2 [d2_stages:0];
  reg [e_len-1:0]  ee  [e_stages:0];



  genvar i;

  // make all inputs signed
  always @(*) aa[a_stages] = signd_a ? a : {1'b0, a}; //spyglass disable W164a W164b
  always @(*) bb[b_stages] = signd_b ? b : {1'b0, b}; //spyglass disable W164a W164b
  generate if (width_b2>0) begin
    (* keep ="true" *) reg [b2_len-1:0] b2_keep;
    always @(*) b2_keep = signd_b2 ? b2 : {1'b0, b2}; //spyglass disable W164a W164b
    always @(*) bb2[b2_stages] = b2_keep;
  end endgenerate
  always @(*) cc[c_stages] = signd_c ? c : {1'b0, c}; //spyglass disable W164a W164b
  always @(*) dd[d_stages] = signd_d ? d : {1'b0, d}; //spyglass disable W164a W164b
  generate if (width_d2>0) begin
    (* keep ="true" *) reg [d2_len-1:0] d2_keep;
    always @(*) d2_keep = signd_d2 ? d2 : {1'b0, d2}; //spyglass disable W164a W164b
    always @(*) dd2[d2_stages] = d2_keep;
  end endgenerate

  generate if (use_const>0) begin
    always @(*) ee[e_stages] = signd_e ? cst : {1'b0, cst}; //spyglass disable W164a W164b

    // input registers
    if (e_stages>0) begin
    for(i = e_stages-1; i >= 0; i=i-1) begin:in_pipe_e
      if (clock_edge == 1'b1) begin:pos
        always @(posedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
      end else begin:neg
        always @(negedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
      end
    end end
  end endgenerate
  generate if (a_stages>0) begin
  for(i = a_stages-1; i >= 0; i=i-1) begin:in_pipe_a
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (b_stages>0) begin
  for(i = b_stages-1; i >= 0; i=i-1) begin:in_pipe_b
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];
    end
  end end endgenerate
  generate if (c_stages>0) begin
  for(i = c_stages-1; i >= 0; i=i-1) begin:in_pipe_c
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (d_stages>0) begin
  for(i = d_stages-1; i >= 0; i=i-1) begin:in_pipe_d
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) dd[i] <= dd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) dd[i] <= dd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (b2_stages>0) begin
  for(i = b2_stages-1; i >= 0; i=i-1) begin:in_pipe_b2
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb2[i] <= bb2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb2[i] <= bb2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (d2_stages>0) begin
  for(i = d2_stages-1; i >= 0; i=i-1) begin:in_pipe_d2
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) dd2[i] <= dd2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) dd2[i] <= dd2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg [bb2_len-1:0] b_bb2[preadd_ab_stages:0];
  reg [dd2_len-1:0] d_dd2[preadd_cd_stages:0];

  //perform first preadd
  generate
    if (width_b2>0) begin
      if (add_b2) begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]) + $signed(bb2[0]); end
      else        begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]) - $signed(bb2[0]); end
    end else      begin always @(*) b_bb2[preadd_ab_stages] = $signed(bb[0]); end
  endgenerate
  generate if (preadd_ab_stages>0) begin
  for(i = preadd_ab_stages-1; i >= 0; i=i-1) begin:preaddab_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) b_bb2[i] <= b_bb2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) b_bb2[i] <= b_bb2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  //perform second preadd
  generate
    if (width_d2>0) begin
      if (add_d2) begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]) + $signed(dd2[0]); end
      else        begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]) - $signed(dd2[0]); end
    end else      begin always @(*) d_dd2[preadd_cd_stages] = $signed(dd[0]); end
  endgenerate
  generate if (preadd_cd_stages>0) begin
  for(i = preadd_cd_stages-1; i >= 0; i=i-1) begin:preaddcd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) d_dd2[i] <= d_dd2[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) d_dd2[i] <= d_dd2[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // perform first multiplication
  reg [axb_len-1:0] axb[axb_stages:0];

  always @(*) axb[axb_stages] = $signed(aa[0]) * $signed(b_bb2[0]);
  generate if (axb_stages>0) begin
  for(i = axb_stages-1; i >= 0; i=i-1) begin:axb_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];
    end
  end end endgenerate

  // perform second multiplication
  reg [cxd_len-1:0] cxd[cxd_stages:0];

  always @(*) cxd[cxd_stages] = $signed(cc[0]) * $signed(d_dd2[0]);
  generate if (cxd_stages>0) begin
  for(i = cxd_stages-1; i >= 0; i=i-1) begin:cxd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cxd[i] <= cxd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cxd[i] <= cxd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg [z_len-1:0]  zz[stages-1:0];
  generate
    if (use_const>1) begin
      reg [z_len-1:0] aux_val;
      if ( isadd) begin
        always @(*) aux_val = $signed(axb[0]) + $signed(cxd[0]);
      end else begin
        always @(*) aux_val = $signed(axb[0]) - $signed(cxd[0]);
      end
      always @(*) zz[stages-1] = $signed(ee[0]) + $signed(aux_val) ;
    end else begin
      if (use_const>0) begin
        if ( isadd) begin always @(*) zz[stages-1] = $signed(axb[0]) + $signed(cxd[0]) + $signed(ee[0]); end else
                    begin always @(*) zz[stages-1] = $signed(axb[0]) - $signed(cxd[0]) + $signed(ee[0]); end
      end else begin
        if ( isadd) begin always @(*) zz[stages-1] = $signed(axb[0]) + $signed(cxd[0]); end else
                    begin always @(*) zz[stages-1] = $signed(axb[0]) - $signed(cxd[0]); end
      end
    end
  endgenerate

  // Output registers:
  generate if (stages>1) begin
  for(i = stages-2; i >= 0; i=i-1) begin:out_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // adjust output
  assign z = zz[0];
endmodule // mgc_mul2add1_pipe

//------> /cad/mentor/2024.2_1/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)
// suppress_sim_read_addr_range_errs:  0 - report errors  1 - suppress errors

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 ,
  parameter suppress_sim_read_addr_range_errs = 1 
  
)( clk,clken,d,q,radr,re,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input  re;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" , syn_ramstyle = "block" *)
  reg [data_width-1:0] mem [depth-1:0];
  integer j;
  initial for (j = 0; j < depth; j = j + 1) mem[j] = 0;
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr READ_ENABLE re
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg re_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
          re_reg <= re;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./PECore.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   grgriff@iron-03
//  Generated date: Tue Jan 20 01:47:23 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_PECoreRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_PECoreRun_fsm (
  clk, rst, PECoreRun_wen, fsm_output
);
  input clk;
  input rst;
  input PECoreRun_wen;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for PECore_PECore_PECoreRun_PECoreRun_fsm_1
  parameter
    PECoreRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : PECore_PECore_PECoreRun_PECoreRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // PECoreRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= PECoreRun_rlp_C_0;
    end
    else if ( PECoreRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_staller
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_staller (
  clk, rst, PECoreRun_wen, PECoreRun_wten, act_port_Push_mioi_wen_comp, rva_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PECoreRun_wen;
  output PECoreRun_wten;
  input act_port_Push_mioi_wen_comp;
  input rva_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg PECoreRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign PECoreRun_wen = act_port_Push_mioi_wen_comp & rva_out_Push_mioi_wen_comp;
  assign PECoreRun_wten = PECoreRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECoreRun_wten_reg <= 1'b0;
    end
    else begin
      PECoreRun_wten_reg <= ~ PECoreRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_wait_dp (
  weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      Datapath_for_4_ProductSum_for_acc_5_cmp_en, Datapath_for_4_ProductSum_for_acc_5_cmp_21_en,
      PECoreRun_wen, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo, weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg,
      Datapath_for_4_ProductSum_for_acc_5_cmp_cgo, Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg,
      Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_21, Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg_21
);
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output Datapath_for_4_ProductSum_for_acc_5_cmp_en;
  output Datapath_for_4_ProductSum_for_acc_5_cmp_21_en;
  input PECoreRun_wen;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg;
  input Datapath_for_4_ProductSum_for_acc_5_cmp_cgo;
  input Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg;
  input Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_21;
  input Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg_21;



  // Interconnect Declarations for Component Instantiations 
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_en = ~(PECoreRun_wen & (Datapath_for_4_ProductSum_for_acc_5_cmp_cgo
      | Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg));
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_21_en = ~(PECoreRun_wen & (Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_21
      | Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg_21));
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  PECoreRun_wen, rva_out_Push_mioi_oswt, rva_out_Push_mioi_biwt, rva_out_Push_mioi_bdwt,
      rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & PECoreRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt)
      & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & rva_out_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt,
      start_PopNB_mioi_biwt_pff, start_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_biwt_pff;
  input start_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & PECoreRun_wen;
  assign start_PopNB_mioi_biwt = (~ PECoreRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_biwt_pff = PECoreRun_wen & start_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp (
  clk, rst, act_port_Push_mioi_oswt, act_port_Push_mioi_wen_comp, act_port_Push_mioi_biwt,
      act_port_Push_mioi_bdwt, act_port_Push_mioi_bcwt, act_port_Push_mioi_m_data_rsc_dat,
      act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff
);
  input clk;
  input rst;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input act_port_Push_mioi_biwt;
  input act_port_Push_mioi_bdwt;
  output act_port_Push_mioi_bcwt;
  reg act_port_Push_mioi_bcwt;
  output [255:0] act_port_Push_mioi_m_data_rsc_dat;
  input [255:0] act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_wen_comp = (~ act_port_Push_mioi_oswt) | act_port_Push_mioi_biwt
      | act_port_Push_mioi_bcwt;
  assign act_port_Push_mioi_m_data_rsc_dat = {16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[239:224])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[207:192])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[175:160])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[143:128])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[111:96])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[79:64])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[47:32])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[15:0])};
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_Push_mioi_bcwt <= ~((~(act_port_Push_mioi_bcwt | act_port_Push_mioi_biwt))
          | act_port_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl (
  PECoreRun_wen, act_port_Push_mioi_oswt, act_port_Push_mioi_biwt, act_port_Push_mioi_bdwt,
      act_port_Push_mioi_bcwt, act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      act_port_Push_mioi_ccs_ccore_done_sync_vld, act_port_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_biwt;
  output act_port_Push_mioi_bdwt;
  input act_port_Push_mioi_bcwt;
  output act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input act_port_Push_mioi_ccs_ccore_done_sync_vld;
  input act_port_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_bdwt = act_port_Push_mioi_oswt & PECoreRun_wen;
  assign act_port_Push_mioi_biwt = act_port_Push_mioi_oswt & (~ act_port_Push_mioi_bcwt)
      & act_port_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & act_port_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
    (
  clk, rst, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt,
      input_port_PopNB_mioi_return_rsc_z_mxwt, input_port_PopNB_mioi_biwt, input_port_PopNB_mioi_bdwt,
      input_port_PopNB_mioi_data_data_data_rsc_z, input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [63:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_biwt;
  input input_port_PopNB_mioi_bdwt;
  input [63:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  input [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  input input_port_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg input_port_PopNB_mioi_bcwt;
  reg [63:0] input_port_PopNB_mioi_data_data_data_rsc_z_bfwt;
  reg [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt;
  reg input_port_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_data_data_data_rsc_z_mxwt = MUX_v_64_2_2(input_port_PopNB_mioi_data_data_data_rsc_z,
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt = MUX_v_8_2_2(input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z,
      input_port_PopNB_mioi_return_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      input_port_PopNB_mioi_bcwt <= ~((~(input_port_PopNB_mioi_bcwt | input_port_PopNB_mioi_biwt))
          | input_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= 8'b00000000;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( input_port_PopNB_mioi_biwt ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= input_port_PopNB_mioi_data_data_data_rsc_z;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= input_port_PopNB_mioi_data_logical_addr_rsc_z;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= input_port_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
    (
  PECoreRun_wen, PECoreRun_wten, input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_biwt,
      input_port_PopNB_mioi_bdwt, input_port_PopNB_mioi_biwt_pff, input_port_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output input_port_PopNB_mioi_biwt;
  output input_port_PopNB_mioi_bdwt;
  output input_port_PopNB_mioi_biwt_pff;
  input input_port_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_bdwt = input_port_PopNB_mioi_oswt & PECoreRun_wen;
  assign input_port_PopNB_mioi_biwt = (~ PECoreRun_wten) & input_port_PopNB_mioi_oswt;
  assign input_port_PopNB_mioi_biwt_pff = PECoreRun_wen & input_port_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [63:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [63:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [63:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  reg [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_64_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_20_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4, rva_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= 20'b00000000000000000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & PECoreRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ PECoreRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = PECoreRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, PECoreRun_wen, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_PECoreRun, rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [63:0] rva_out_dat;
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [63:0] rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_oswt_pff(rva_out_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi (
  clk, rst, start_vld, start_rdy, start_dat, PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_vld(start_vld),
      .this_rdy(start_rdy),
      .this_dat(start_dat),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_biwt_pff(start_PopNB_mioi_biwt_iff),
      .start_PopNB_mioi_oswt_pff(start_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi (
  clk, rst, act_port_vld, act_port_rdy, act_port_dat, PECoreRun_wen, act_port_Push_mioi_oswt,
      act_port_Push_mioi_wen_comp, act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff,
      act_port_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input [255:0] act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff;
  input act_port_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_port_Push_mioi_biwt;
  wire act_port_Push_mioi_bdwt;
  wire act_port_Push_mioi_bcwt;
  wire [255:0] act_port_Push_mioi_m_data_rsc_dat;
  wire act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire act_port_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [255:0] nl_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff;
  assign nl_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff
      = {16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[239:224])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[207:192])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[175:160])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[143:128])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[111:96])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[79:64])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[47:32])
      , 16'b0000000000000000 , (act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[15:0])};
  PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push  act_port_Push_mioi
      (
      .this_vld(act_port_vld),
      .this_rdy(act_port_rdy),
      .this_dat(act_port_dat),
      .m_data_rsc_dat(act_port_Push_mioi_m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt),
      .act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .act_port_Push_mioi_ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .act_port_Push_mioi_oswt_pff(act_port_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt),
      .act_port_Push_mioi_m_data_rsc_dat(act_port_Push_mioi_m_data_rsc_dat),
      .act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff(nl_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[255:0])
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi (
  clk, rst, input_port_vld, input_port_rdy, input_port_dat, PECoreRun_wen, PECoreRun_wten,
      input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt, input_port_PopNB_mioi_return_rsc_z_mxwt,
      input_port_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input input_port_vld;
  output input_port_rdy;
  input [73:0] input_port_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output [63:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_port_PopNB_mioi_biwt;
  wire input_port_PopNB_mioi_bdwt;
  wire [63:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  wire input_port_PopNB_mioi_return_rsc_z;
  wire input_port_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB  input_port_PopNB_mioi
      (
      .this_vld(input_port_vld),
      .this_rdy(input_port_rdy),
      .this_dat(input_port_dat),
      .data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .return_rsc_z(input_port_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(input_port_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(input_port_PopNB_mioi_oswt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_biwt_pff(input_port_PopNB_mioi_biwt_iff),
      .input_port_PopNB_mioi_oswt_pff(input_port_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .input_port_PopNB_mioi_return_rsc_z(input_port_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt,
      rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [96:0] rva_in_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [63:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [63:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG, weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d, Datapath_for_4_ProductSum_for_acc_5_cmp_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_c, Datapath_for_4_ProductSum_for_acc_5_cmp_en,
      Datapath_for_4_ProductSum_for_acc_5_cmp_z, Datapath_for_4_ProductSum_for_acc_5_cmp_1_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_1_c, Datapath_for_4_ProductSum_for_acc_5_cmp_1_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_2_a, Datapath_for_4_ProductSum_for_acc_5_cmp_2_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_2_z, Datapath_for_4_ProductSum_for_acc_5_cmp_3_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_3_c, Datapath_for_4_ProductSum_for_acc_5_cmp_3_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_4_a, Datapath_for_4_ProductSum_for_acc_5_cmp_4_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_4_z, Datapath_for_4_ProductSum_for_acc_5_cmp_5_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_5_c, Datapath_for_4_ProductSum_for_acc_5_cmp_5_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_a, Datapath_for_4_ProductSum_for_acc_5_cmp_6_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_z, Datapath_for_4_ProductSum_for_acc_5_cmp_7_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_7_c, Datapath_for_4_ProductSum_for_acc_5_cmp_7_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_8_a, Datapath_for_4_ProductSum_for_acc_5_cmp_8_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_8_z, Datapath_for_4_ProductSum_for_acc_5_cmp_9_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_9_c, Datapath_for_4_ProductSum_for_acc_5_cmp_9_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_10_a, Datapath_for_4_ProductSum_for_acc_5_cmp_10_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_10_z, Datapath_for_4_ProductSum_for_acc_5_cmp_11_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_11_c, Datapath_for_4_ProductSum_for_acc_5_cmp_11_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_12_a, Datapath_for_4_ProductSum_for_acc_5_cmp_12_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_12_z, Datapath_for_4_ProductSum_for_acc_5_cmp_13_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_13_c, Datapath_for_4_ProductSum_for_acc_5_cmp_13_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_14_a, Datapath_for_4_ProductSum_for_acc_5_cmp_14_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_14_z, Datapath_for_4_ProductSum_for_acc_5_cmp_15_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_15_c, Datapath_for_4_ProductSum_for_acc_5_cmp_15_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_16_a, Datapath_for_4_ProductSum_for_acc_5_cmp_16_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_16_z, Datapath_for_4_ProductSum_for_acc_5_cmp_17_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_17_c, Datapath_for_4_ProductSum_for_acc_5_cmp_17_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_18_a, Datapath_for_4_ProductSum_for_acc_5_cmp_18_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_18_z, Datapath_for_4_ProductSum_for_acc_5_cmp_19_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_19_c, Datapath_for_4_ProductSum_for_acc_5_cmp_19_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_20_a, Datapath_for_4_ProductSum_for_acc_5_cmp_20_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_20_z, Datapath_for_4_ProductSum_for_acc_5_cmp_21_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_21_b, Datapath_for_4_ProductSum_for_acc_5_cmp_21_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_21_d, Datapath_for_4_ProductSum_for_acc_5_cmp_21_en,
      Datapath_for_4_ProductSum_for_acc_5_cmp_21_z, Datapath_for_4_ProductSum_for_acc_5_cmp_22_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_22_c, Datapath_for_4_ProductSum_for_acc_5_cmp_22_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_23_a, Datapath_for_4_ProductSum_for_acc_5_cmp_23_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_23_z, Datapath_for_4_ProductSum_for_acc_5_cmp_24_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_24_c, Datapath_for_4_ProductSum_for_acc_5_cmp_24_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_25_a, Datapath_for_4_ProductSum_for_acc_5_cmp_25_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_25_z, Datapath_for_4_ProductSum_for_acc_5_cmp_26_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_26_c, Datapath_for_4_ProductSum_for_acc_5_cmp_26_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_27_a, Datapath_for_4_ProductSum_for_acc_5_cmp_27_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_27_z, Datapath_for_4_ProductSum_for_acc_5_cmp_28_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_28_c, Datapath_for_4_ProductSum_for_acc_5_cmp_28_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_29_a, Datapath_for_4_ProductSum_for_acc_5_cmp_29_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_29_z, Datapath_for_4_ProductSum_for_acc_5_cmp_30_a,
      Datapath_for_4_ProductSum_for_acc_5_cmp_30_c, Datapath_for_4_ProductSum_for_acc_5_cmp_30_z,
      Datapath_for_4_ProductSum_for_acc_5_cmp_31_a, Datapath_for_4_ProductSum_for_acc_5_cmp_31_c,
      Datapath_for_4_ProductSum_for_acc_5_cmp_31_z, Datapath_for_4_ProductSum_for_acc_5_cmp_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_pff, Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_pff,
      Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff, weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [73:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [96:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [63:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_c;
  output Datapath_for_4_ProductSum_for_acc_5_cmp_en;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_b;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_c;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_d;
  output Datapath_for_4_ProductSum_for_acc_5_cmp_21_en;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_a;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_c;
  input [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_z;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_pff;
  output [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff;


  // Interconnect Declarations
  wire PECoreRun_wen;
  wire PECoreRun_wten;
  wire [63:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [63:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  wire input_port_PopNB_mioi_return_rsc_z_mxwt;
  wire act_port_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
  wire fsm_output;
  wire pe_config_UpdateManagerCounter_if_if_unequal_tmp;
  wire [7:0] weight_mem_write_arbxbar_xbar_for_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_7_false_1_operator_7_false_1_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_1_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp;
  wire while_mux_1304_tmp;
  wire while_mux_1303_tmp;
  wire while_mux_1302_tmp;
  wire while_mux_1301_tmp;
  wire while_mux_1300_tmp;
  wire while_mux_1299_tmp;
  wire while_mux_1297_tmp;
  wire while_mux_1296_tmp;
  wire while_mux_1295_tmp;
  wire while_mux_1294_tmp;
  wire while_mux_1293_tmp;
  wire while_mux_1292_tmp;
  wire while_mux_1291_tmp;
  wire while_mux_1290_tmp;
  wire while_mux_1289_tmp;
  wire while_mux_1288_tmp;
  wire while_mux_1287_tmp;
  wire while_mux_1286_tmp;
  wire while_mux_1285_tmp;
  wire while_mux_1284_tmp;
  wire while_mux_1276_tmp;
  wire while_mux_1275_tmp;
  wire while_mux_1274_tmp;
  wire while_mux_1273_tmp;
  wire while_mux_1272_tmp;
  wire while_mux_1271_tmp;
  wire while_mux_1270_tmp;
  wire while_mux_1254_tmp;
  wire while_mux_1251_tmp;
  wire while_mux_1250_tmp;
  wire while_mux_1249_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_103_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_99_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_75_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_23_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_1_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_111_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  wire and_dcpl_4;
  wire and_dcpl_5;
  wire and_dcpl_6;
  wire and_dcpl_22;
  wire and_dcpl_25;
  wire and_dcpl_27;
  wire and_dcpl_28;
  wire and_dcpl_30;
  wire mux_tmp;
  wire or_tmp;
  wire and_dcpl_43;
  wire and_dcpl_44;
  wire or_tmp_2;
  wire not_tmp_33;
  wire or_tmp_60;
  wire and_dcpl_74;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_87;
  wire and_dcpl_89;
  wire and_dcpl_90;
  wire or_dcpl_59;
  wire or_dcpl_68;
  wire and_dcpl_140;
  wire and_dcpl_141;
  wire and_dcpl_142;
  wire and_dcpl_143;
  wire and_dcpl_144;
  wire and_dcpl_145;
  wire and_dcpl_146;
  wire and_dcpl_147;
  wire and_dcpl_153;
  wire and_dcpl_158;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_173;
  wire and_dcpl_174;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_179;
  wire and_dcpl_180;
  wire and_dcpl_182;
  wire and_dcpl_183;
  wire and_dcpl_185;
  wire and_dcpl_186;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_194;
  wire and_dcpl_198;
  wire and_dcpl_201;
  wire or_dcpl_135;
  wire or_dcpl_141;
  wire and_dcpl_203;
  wire and_dcpl_206;
  wire and_dcpl_207;
  wire and_dcpl_208;
  wire and_dcpl_209;
  wire and_dcpl_211;
  wire or_tmp_84;
  wire mux_tmp_60;
  wire mux_tmp_62;
  wire or_tmp_94;
  wire or_tmp_95;
  wire and_dcpl_240;
  wire and_dcpl_244;
  wire and_dcpl_245;
  wire and_dcpl_248;
  wire and_dcpl_267;
  wire or_tmp_111;
  wire and_dcpl_284;
  wire and_dcpl_297;
  wire and_dcpl_305;
  wire and_dcpl_308;
  wire and_dcpl_309;
  wire not_tmp_182;
  wire and_dcpl_325;
  wire and_dcpl_337;
  wire and_dcpl_349;
  wire and_dcpl_350;
  wire and_dcpl_357;
  wire and_dcpl_375;
  wire and_dcpl_393;
  wire and_dcpl_406;
  wire and_dcpl_417;
  wire and_dcpl_434;
  wire and_dcpl_435;
  wire mux_tmp_97;
  wire and_dcpl_441;
  wire and_dcpl_476;
  wire and_dcpl_480;
  wire and_dcpl_486;
  wire mux_tmp_98;
  wire mux_tmp_99;
  wire and_dcpl_489;
  wire mux_tmp_102;
  wire mux_tmp_103;
  wire not_tmp_264;
  wire not_tmp_267;
  wire not_tmp_270;
  wire or_tmp_164;
  wire nor_tmp_47;
  wire mux_tmp_113;
  wire not_tmp_274;
  wire not_tmp_277;
  wire or_tmp_178;
  wire nor_tmp_50;
  wire mux_tmp_123;
  wire not_tmp_281;
  wire or_dcpl_218;
  wire and_dcpl_543;
  wire and_dcpl_544;
  wire and_dcpl_545;
  wire or_dcpl_227;
  wire or_dcpl_228;
  wire or_dcpl_239;
  wire or_dcpl_240;
  wire and_dcpl_594;
  wire and_dcpl_595;
  wire and_dcpl_596;
  wire and_dcpl_597;
  wire and_dcpl_599;
  wire and_dcpl_603;
  wire or_dcpl_275;
  wire or_dcpl_278;
  wire or_dcpl_283;
  wire nor_tmp_58;
  wire or_tmp_206;
  wire mux_tmp_152;
  wire or_tmp_208;
  wire or_tmp_209;
  wire mux_tmp_153;
  wire not_tmp_425;
  wire or_tmp_223;
  wire or_tmp_229;
  wire and_dcpl_632;
  wire or_tmp_243;
  wire or_tmp_245;
  wire mux_tmp_178;
  wire or_tmp_247;
  wire or_tmp_249;
  wire or_tmp_250;
  wire or_tmp_252;
  wire or_tmp_254;
  wire or_tmp_259;
  wire or_tmp_262;
  wire mux_tmp_197;
  wire or_tmp_266;
  wire nor_tmp_117;
  wire or_tmp_272;
  wire nor_tmp_120;
  wire or_tmp_278;
  wire and_dcpl_634;
  wire or_tmp_287;
  wire or_tmp_292;
  wire or_tmp_294;
  wire or_tmp_296;
  wire mux_tmp_220;
  wire or_tmp_300;
  wire or_tmp_303;
  wire or_tmp_304;
  wire mux_tmp_236;
  wire or_tmp_305;
  wire or_tmp_306;
  wire or_tmp_308;
  wire nor_tmp_154;
  wire or_tmp_310;
  wire or_tmp_311;
  wire or_tmp_312;
  wire or_tmp_314;
  wire mux_tmp_237;
  wire mux_tmp_239;
  wire and_dcpl_637;
  wire mux_tmp_252;
  wire and_dcpl_639;
  wire and_dcpl_642;
  wire and_dcpl_643;
  wire and_dcpl_644;
  wire or_tmp_327;
  wire or_tmp_329;
  wire mux_tmp_255;
  wire mux_tmp_258;
  wire mux_tmp_261;
  wire or_tmp_334;
  wire or_tmp_339;
  wire or_tmp_342;
  wire or_tmp_347;
  wire nor_tmp_181;
  wire or_tmp_353;
  wire nor_tmp_184;
  wire or_tmp_359;
  wire and_dcpl_647;
  wire or_tmp_368;
  wire or_tmp_373;
  wire or_tmp_375;
  wire or_tmp_377;
  wire mux_tmp_290;
  wire or_tmp_379;
  wire or_tmp_383;
  wire or_tmp_388;
  wire or_tmp_391;
  wire or_tmp_392;
  wire or_tmp_393;
  wire or_tmp_396;
  wire or_tmp_397;
  wire or_tmp_398;
  wire mux_tmp_296;
  wire mux_tmp_297;
  wire and_dcpl_648;
  wire and_dcpl_652;
  wire and_dcpl_655;
  wire and_dcpl_656;
  wire and_dcpl_657;
  wire and_dcpl_661;
  wire and_dcpl_662;
  wire and_dcpl_665;
  wire or_dcpl_296;
  wire while_and_24_cse;
  wire [3:0] pe_config_manager_counter_sva_mx1;
  wire [4:0] operator_4_false_acc_sdt_sva_1;
  wire [5:0] nl_operator_4_false_acc_sdt_sva_1;
  reg [3:0] pe_config_num_manager_sva;
  wire state_0_sva_mx1;
  wire while_if_and_tmp_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiWrite_switch_lp_nor_tmp_1;
  reg pe_config_is_valid_sva;
  reg pe_config_is_zero_first_sva;
  reg pe_manager_zero_active_sva;
  reg pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  reg pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  reg PECore_UpdateFSM_switch_lp_and_7_itm_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
  reg PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  reg [8:0] operator_8_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_8_false_acc_sdt_sva_1;
  wire PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  wire PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1;
  reg PECore_RunFSM_switch_lp_nor_tmp_1;
  reg [1:0] state_2_1_sva;
  reg state_0_sva;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  wire nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_5_mux_2_mx0w3;
  wire nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_4_mux_2_mx0w2;
  wire weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  reg Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1;
  reg PECore_RunFSM_switch_lp_equal_tmp_1_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  reg weight_mem_run_3_for_land_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg input_read_req_valid_lpi_1_dfm_1_10;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8;
  reg rva_in_reg_rw_sva_10;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_10;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  wire PECore_UpdateFSM_switch_lp_equal_tmp_6;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  wire PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
  wire PECore_UpdateFSM_switch_lp_nor_tmp_1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
  wire [7:0] pe_config_input_counter_sva_mx1;
  wire [8:0] operator_16_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_16_false_acc_sdt_sva_1;
  reg [7:0] pe_manager_num_input_sva;
  reg [7:0] pe_config_num_output_sva;
  wire PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10;
  reg weight_mem_run_3_for_land_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  wire PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  reg PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
  wire weight_mem_run_3_for_land_lpi_1_dfm_1_1;
  wire weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  wire weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  wire weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_1_itm_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  wire weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_127_sva_1;
  reg input_write_req_valid_lpi_1_dfm_1_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1;
  wire input_write_req_valid_lpi_1_dfm_5;
  wire input_mem_banks_write_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1;
  reg [14:0] pe_manager_base_input_sva;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1;
  reg rva_in_reg_rw_sva_5;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_4;
  wire PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3;
  reg rva_in_reg_rw_sva_st_1_10;
  reg rva_in_reg_rw_sva_9;
  reg input_read_req_valid_lpi_1_dfm_1_9;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
  reg rva_in_reg_rw_sva_st_1_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
  reg while_stage_0_11;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  reg rva_in_reg_rw_sva_st_1_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  reg while_stage_0_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
  reg rva_in_reg_rw_sva_st_1_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1;
  reg while_stage_0_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
  reg rva_in_reg_rw_sva_4;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5;
  reg weight_mem_read_arbxbar_arbiters_next_7_6_sva;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  reg while_stage_0_4;
  reg weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  reg while_stage_0_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2;
  reg rva_in_reg_rw_sva_st_1_4;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
  reg while_stage_0_3;
  reg PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  reg [1:0] state_2_1_sva_dfm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
  reg rva_in_reg_rw_sva_st_1_3;
  reg rva_in_reg_rw_sva_st_1_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  reg input_read_req_valid_lpi_1_dfm_1_8;
  reg rva_in_reg_rw_sva_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
  reg while_stage_0_10;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
  reg rva_in_reg_rw_sva_st_1_7;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  reg input_read_req_valid_lpi_1_dfm_1_7;
  reg rva_in_reg_rw_sva_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
  reg while_stage_0_9;
  reg input_read_req_valid_lpi_1_dfm_1_2;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
  reg input_read_req_valid_lpi_1_dfm_1_6;
  reg rva_in_reg_rw_sva_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
  reg input_read_req_valid_lpi_1_dfm_1_1;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
  reg rva_in_reg_rw_sva_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2;
  reg input_read_req_valid_lpi_1_dfm_1_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1;
  reg [3:0] while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
  reg while_stage_0_8;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3;
  reg weight_mem_run_3_for_5_and_132_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10;
  reg while_stage_0_12;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_9;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_9;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_2;
  reg while_and_1126_itm_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
  reg weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_2_sva;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs;
  wire operator_7_false_1_operator_7_false_1_or_mdf_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1;
  wire operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_3_2_0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_2_2_0;
  reg [14:0] weight_read_addrs_7_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_5_lpi_1_dfm_1;
  reg [14:0] pe_manager_base_weight_sva;
  reg [14:0] weight_read_addrs_3_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_1_lpi_1_dfm_1;
  wire [14:0] pe_manager_base_weight_sva_mx2;
  wire [3:0] pe_manager_base_weight_sva_mx1_3_0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  wire [11:0] nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_2;
  reg [7:0] while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4;
  wire [7:0] input_write_addrs_lpi_1_dfm_2;
  wire PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
  wire weight_mem_banks_read_1_for_mux_cse;
  wire weight_mem_banks_read_1_for_mux_1_cse;
  wire weight_mem_banks_read_1_for_mux_4_cse;
  wire weight_mem_banks_read_1_for_mux_5_cse;
  wire weight_mem_banks_read_1_for_mux_8_cse;
  wire weight_mem_banks_read_1_for_mux_9_cse;
  wire weight_mem_banks_read_1_for_mux_12_cse;
  wire weight_mem_banks_read_1_for_mux_13_cse;
  wire weight_mem_banks_read_1_for_mux_16_cse;
  wire weight_mem_banks_read_1_for_mux_17_cse;
  wire weight_mem_banks_read_1_for_mux_20_cse;
  wire weight_mem_banks_read_1_for_mux_21_cse;
  wire weight_mem_banks_read_1_for_mux_24_cse;
  wire weight_mem_banks_read_1_for_mux_25_cse;
  wire weight_mem_banks_read_1_for_mux_28_cse;
  wire weight_mem_banks_read_1_for_mux_29_cse;
  wire weight_mem_banks_write_if_for_if_mux_8_cse;
  wire weight_mem_banks_write_if_for_if_mux_9_cse;
  wire weight_mem_banks_read_for_mux_cse;
  wire weight_mem_banks_read_for_mux_1_cse;
  wire weight_mem_banks_write_if_for_if_mux_12_cse;
  wire weight_mem_banks_write_if_for_if_mux_13_cse;
  wire weight_mem_banks_read_for_mux_4_cse;
  wire weight_mem_banks_read_for_mux_5_cse;
  wire weight_mem_banks_write_if_for_if_mux_16_cse;
  wire weight_mem_banks_write_if_for_if_mux_17_cse;
  wire weight_mem_banks_read_for_mux_8_cse;
  wire weight_mem_banks_read_for_mux_9_cse;
  wire weight_mem_banks_write_if_for_if_mux_20_cse;
  wire weight_mem_banks_write_if_for_if_mux_21_cse;
  wire weight_mem_banks_read_for_mux_12_cse;
  wire weight_mem_banks_read_for_mux_13_cse;
  wire weight_mem_banks_write_if_for_if_mux_24_cse;
  wire weight_mem_banks_write_if_for_if_mux_25_cse;
  wire weight_mem_banks_read_for_mux_16_cse;
  wire weight_mem_banks_read_for_mux_17_cse;
  wire weight_mem_banks_write_if_for_if_mux_28_cse;
  wire weight_mem_banks_write_if_for_if_mux_29_cse;
  wire weight_mem_banks_read_for_mux_20_cse;
  wire weight_mem_banks_read_for_mux_21_cse;
  wire weight_mem_banks_write_if_for_if_mux_32_cse;
  wire weight_mem_banks_write_if_for_if_mux_33_cse;
  wire weight_mem_banks_read_for_mux_24_cse;
  wire weight_mem_banks_read_for_mux_25_cse;
  wire weight_mem_banks_write_if_for_if_mux_36_cse;
  wire weight_mem_banks_write_if_for_if_mux_37_cse;
  wire weight_mem_banks_read_for_mux_28_cse;
  wire weight_mem_banks_read_for_mux_29_cse;
  wire input_mem_banks_write_1_if_for_if_mux_cse;
  wire input_mem_banks_write_1_if_for_if_mux_1_cse;
  wire input_mem_banks_read_1_for_mux_cse;
  wire input_mem_banks_read_1_for_mux_1_cse;
  wire input_mem_banks_write_if_for_if_mux_cse;
  wire input_mem_banks_write_if_for_if_mux_1_cse;
  wire input_mem_banks_read_for_mux_cse;
  wire input_mem_banks_read_for_mux_1_cse;
  reg reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_31_cse;
  reg reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_21_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_act_port_Push_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire rva_out_reg_data_and_cse;
  wire weight_port_read_out_data_and_10_cse;
  wire weight_port_read_out_data_and_18_cse;
  wire weight_port_read_out_data_and_24_cse;
  wire weight_port_read_out_data_and_32_cse;
  wire weight_port_read_out_data_and_56_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_cse;
  reg reg_rva_in_reg_rw_sva_st_1_1_cse;
  wire or_220_cse;
  reg [2:0] reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse;
  wire operator_15_false_1_and_cse;
  wire pe_config_num_manager_and_cse;
  wire PECore_DecodeAxiWrite_switch_lp_and_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
  wire or_296_cse;
  wire or_261_cse;
  wire or_286_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_cse;
  reg reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
  wire pe_manager_num_input_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_56_cse;
  wire Arbiter_8U_Roundrobin_pick_and_36_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_44_cse;
  wire Arbiter_8U_Roundrobin_pick_and_30_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_32_cse;
  wire Arbiter_8U_Roundrobin_pick_and_24_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_20_cse;
  wire Arbiter_8U_Roundrobin_pick_and_18_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_8_cse;
  wire Arbiter_8U_Roundrobin_pick_and_12_cse;
  wire [1:0] state_mux_1_cse;
  wire and_301_cse;
  wire and_713_cse;
  wire and_715_cse;
  wire and_522_cse;
  wire and_887_cse;
  wire and_889_cse;
  wire and_888_cse;
  wire and_890_cse;
  wire or_38_cse;
  wire and_882_cse;
  wire and_706_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
  wire or_708_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
  wire and_604_cse;
  wire or_231_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  wire while_and_23_cse;
  wire nor_253_cse;
  wire nor_226_cse;
  wire nor_227_cse;
  wire nor_228_cse;
  wire nor_229_cse;
  wire nor_233_cse;
  wire nor_231_cse;
  wire nor_237_cse;
  wire and_121_cse;
  wire nor_242_cse;
  wire nor_246_cse;
  wire nor_260_cse;
  wire nand_31_cse;
  wire and_728_cse;
  wire and_686_cse;
  wire and_679_cse;
  wire and_893_cse;
  wire and_892_cse;
  wire and_891_cse;
  wire and_894_cse;
  wire and_755_cse;
  wire and_756_cse;
  wire and_757_cse;
  wire and_758_cse;
  wire and_761_cse;
  wire and_763_cse;
  wire and_768_cse;
  wire and_772_cse;
  wire and_782_cse;
  wire and_776_cse;
  wire and_781_cse;
  wire and_792_cse;
  wire and_791_cse;
  wire and_794_cse;
  wire and_793_cse;
  wire and_805_cse;
  wire and_804_cse;
  wire and_815_cse;
  wire and_809_cse;
  wire and_820_cse;
  wire and_824_cse;
  wire and_825_cse;
  wire and_822_cse;
  wire and_828_cse;
  wire and_829_cse;
  wire and_826_cse;
  wire and_830_cse;
  wire and_853_cse;
  wire and_854_cse;
  wire and_855_cse;
  wire and_856_cse;
  wire and_859_cse;
  wire and_860_cse;
  wire and_863_cse;
  wire and_864_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse;
  reg Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_4_mx1w0;
  wire operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1;
  wire while_if_and_2_m1c;
  wire mux_142_cse;
  wire pe_config_is_valid_and_cse;
  wire weight_mem_run_3_for_5_and_177_cse;
  wire weight_mem_run_3_for_5_and_197_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_cse;
  wire Arbiter_8U_Roundrobin_pick_and_38_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_69_cse;
  wire Arbiter_8U_Roundrobin_pick_and_50_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_81_cse;
  wire Arbiter_8U_Roundrobin_pick_and_62_cse;
  wire pe_config_input_counter_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse;
  wire PECore_PushAxiRsp_and_2_cse;
  wire and_142_cse;
  wire and_107_cse;
  wire and_114_cse;
  wire and_128_cse;
  wire and_135_cse;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1;
  wire PECore_DecodeAxiWrite_switch_lp_or_5_cse_1;
  wire weight_mem_run_3_for_5_and_175_cse;
  wire weight_mem_run_3_for_5_and_176_cse;
  wire weight_mem_run_3_for_5_and_178_cse;
  wire weight_mem_run_3_for_5_and_182_cse;
  wire weight_mem_run_3_for_5_and_196_cse;
  wire weight_mem_run_3_for_5_and_189_cse;
  wire weight_mem_run_3_for_5_and_203_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_73_cse;
  wire nand_39_cse;
  wire weight_mem_run_3_for_weight_mem_run_3_for_and_4_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0;
  wire and_520_rmff;
  wire and_517_rmff;
  wire and_514_rmff;
  wire and_511_rmff;
  wire and_508_rmff;
  wire and_505_rmff;
  wire and_502_rmff;
  wire and_497_rmff;
  wire and_489_rmff;
  wire and_492_rmff;
  wire and_524_rmff;
  wire and_526_rmff;
  reg [7:0] pe_config_output_counter_sva;
  reg [7:0] pe_config_input_counter_sva;
  reg rva_out_reg_data_63_sva_dfm_4_5;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_5;
  reg rva_out_reg_data_47_sva_dfm_4_5;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_5;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_4;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0;
  reg weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
  reg [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1;
  reg [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1;
  reg [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1;
  reg weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
  reg [63:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
  wire [7:0] weight_port_read_out_data_7_1_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_0_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_3_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_2_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_5_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_4_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_7_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_6_sva_dfm_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
  reg [7:0] weight_port_read_out_data_6_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_6_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_6_3_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_6_2_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_6_5_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_6_4_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_6_7_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_6_6_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_1_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
  reg [7:0] weight_port_read_out_data_1_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
  reg [7:0] weight_port_read_out_data_1_3_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
  reg [7:0] weight_port_read_out_data_1_2_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
  reg [7:0] weight_port_read_out_data_1_5_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004;
  reg [7:0] weight_port_read_out_data_1_4_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005;
  reg [7:0] weight_port_read_out_data_1_7_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_000000;
  reg [7:0] weight_port_read_out_data_1_6_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
  reg [7:0] weight_port_read_out_data_2_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_3_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
  reg [7:0] weight_port_read_out_data_2_2_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
  reg [7:0] weight_port_read_out_data_2_5_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
  reg [7:0] weight_port_read_out_data_2_4_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004;
  reg [7:0] weight_port_read_out_data_2_7_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_sva_1;
  reg [7:0] weight_port_read_out_data_2_6_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005;
  reg [7:0] weight_port_read_out_data_4_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_4_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_4_3_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_4_2_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_4_5_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_4_4_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_4_7_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_4_6_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_port_read_out_data_3_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
  reg [7:0] weight_port_read_out_data_3_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
  reg [7:0] weight_port_read_out_data_3_3_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
  reg [7:0] weight_port_read_out_data_3_2_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
  reg [14:0] weight_write_addrs_lpi_1_dfm_1_2;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_3_2;
  reg [11:0] weight_write_addrs_lpi_1_dfm_1_3_14_3;
  reg [15:0] act_port_reg_data_239_224_sva_dfm_1_2;
  reg [15:0] act_port_reg_data_207_192_sva_dfm_1_2;
  reg [15:0] act_port_reg_data_175_160_sva_dfm_1_2;
  reg [15:0] act_port_reg_data_143_128_sva_dfm_1_2;
  reg [15:0] act_port_reg_data_111_96_sva_dfm_1_2;
  reg [15:0] act_port_reg_data_79_64_sva_dfm_1_1;
  reg [15:0] act_port_reg_data_47_32_sva_dfm_1_2;
  reg [15:0] act_port_reg_data_15_0_sva_dfm_1_2;
  wire or_dcpl_297;
  wire and_dcpl_678;
  wire and_dcpl_679;
  wire or_dcpl_302;
  wire or_dcpl_303;
  reg [63:0] input_mem_banks_read_read_data_lpi_1_dfm_1_4;
  reg [63:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1;
  wire [63:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0;
  wire [55:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_2;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2;
  wire or_713_tmp;
  wire or_718_tmp;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_4;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_2;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_2;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_4;
  wire and_937_cse;
  wire and_938_cse;
  wire and_939_cse;
  wire and_940_cse;
  wire and_941_cse;
  wire and_942_cse;
  wire nor_427_cse;
  wire and_927_cse;
  wire and_928_cse;
  wire and_929_cse;
  wire and_930_cse;
  wire and_931_cse;
  wire and_932_cse;
  wire and_933_cse;
  wire nor_426_cse;
  wire and_536_itm;
  wire nor_413_itm;
  wire [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm;
  wire [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm;
  wire mux_160_itm;
  wire mux_193_itm;
  wire mux_207_itm;
  wire mux_235_itm;
  wire mux_244_itm;
  wire mux_264_itm;
  wire mux_277_itm;
  wire mux_295_itm;
  reg weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_4_sva;
  reg [14:0] pe_manager_base_bias_sva;
  reg pe_config_is_cluster_sva;
  reg pe_config_is_bias_sva;
  reg [3:0] pe_config_manager_counter_sva;
  reg [18:0] accum_vector_data_3_18_0_sva;
  reg [18:0] accum_vector_data_4_18_0_sva;
  reg [18:0] accum_vector_data_2_18_0_sva;
  reg [18:0] accum_vector_data_5_18_0_sva;
  reg [18:0] accum_vector_data_1_18_0_sva;
  reg [18:0] accum_vector_data_6_18_0_sva;
  reg [18:0] accum_vector_data_0_18_0_sva;
  reg [18:0] accum_vector_data_7_18_0_sva;
  reg [15:0] act_port_reg_data_111_96_sva;
  reg [15:0] act_port_reg_data_143_128_sva;
  reg [15:0] act_port_reg_data_79_64_sva;
  reg [15:0] act_port_reg_data_175_160_sva;
  reg [15:0] act_port_reg_data_47_32_sva;
  reg [15:0] act_port_reg_data_207_192_sva;
  reg [15:0] act_port_reg_data_15_0_sva;
  reg [15:0] act_port_reg_data_239_224_sva;
  reg [7:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8;
  reg [63:0] input_mem_banks_bank_a_0_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_1_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_2_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_3_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_4_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_5_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_6_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_7_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_8_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_9_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_10_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_11_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_12_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_13_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_14_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_15_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_16_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_17_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_18_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_19_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_20_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_21_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_22_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_23_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_24_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_25_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_26_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_27_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_28_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_29_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_30_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_31_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_32_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_33_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_34_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_35_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_36_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_37_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_38_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_39_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_40_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_41_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_42_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_43_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_44_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_45_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_46_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_47_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_48_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_49_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_50_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_51_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_52_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_53_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_54_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_55_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_56_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_57_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_58_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_59_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_60_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_61_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_62_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_63_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_64_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_65_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_66_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_67_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_68_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_69_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_70_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_71_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_72_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_73_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_74_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_75_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_76_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_77_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_78_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_79_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_80_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_81_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_82_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_83_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_84_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_85_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_86_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_87_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_88_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_89_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_90_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_91_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_92_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_93_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_94_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_95_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_96_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_97_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_98_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_99_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_100_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_101_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_102_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_103_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_104_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_105_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_106_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_107_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_108_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_109_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_110_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_111_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_112_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_113_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_114_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_115_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_116_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_117_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_118_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_119_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_120_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_121_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_122_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_123_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_124_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_125_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_126_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_127_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_128_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_129_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_130_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_131_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_132_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_133_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_134_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_135_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_136_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_137_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_138_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_139_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_140_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_141_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_142_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_143_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_144_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_145_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_146_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_147_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_148_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_149_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_150_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_151_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_152_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_153_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_154_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_155_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_156_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_157_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_158_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_159_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_160_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_161_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_162_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_163_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_164_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_165_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_166_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_167_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_168_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_169_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_170_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_171_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_172_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_173_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_174_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_175_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_176_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_177_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_178_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_179_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_180_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_181_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_182_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_183_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_184_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_185_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_186_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_187_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_188_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_189_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_190_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_191_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_192_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_193_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_194_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_195_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_196_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_197_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_198_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_199_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_200_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_201_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_202_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_203_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_204_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_205_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_206_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_207_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_208_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_209_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_210_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_211_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_212_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_213_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_214_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_215_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_216_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_217_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_218_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_219_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_220_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_221_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_222_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_223_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_224_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_225_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_226_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_227_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_228_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_229_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_230_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_231_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_232_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_233_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_234_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_235_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_236_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_237_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_238_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_239_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_240_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_241_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_242_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_243_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_244_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_245_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_246_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_247_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_248_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_249_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_250_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_251_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_252_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_253_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_254_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_255_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_2_1_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_1_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_1_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_7_sva_dfm_1;
  reg rva_out_reg_data_24_sva_dfm_6;
  reg rva_out_reg_data_31_sva_dfm_6;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_6;
  reg rva_out_reg_data_16_sva_dfm_6;
  reg rva_out_reg_data_8_sva_dfm_6;
  reg rva_out_reg_data_0_sva_dfm_6;
  reg [63:0] weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1;
  reg [63:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1;
  reg [63:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1;
  reg [63:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_6;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_2;
  reg [7:0] weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2;
  reg [3:0] pe_config_manager_counter_sva_dfm_3_1;
  reg [7:0] input_read_addrs_sva_1_1;
  wire [8:0] nl_input_read_addrs_sva_1_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_2;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_3;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_4;
  reg rva_out_reg_data_63_sva_dfm_4_4;
  reg rva_out_reg_data_47_sva_dfm_4_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_3;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_4;
  reg [63:0] input_mem_banks_read_read_data_sva_1;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_1;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_5;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_1;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_2;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_3;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_4;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_5;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_6;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_7;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_8;
  reg [7:0] pe_config_output_counter_sva_dfm_1;
  reg [7:0] pe_config_input_counter_sva_dfm_1;
  reg [63:0] rva_in_reg_data_sva_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_2;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_1;
  reg [10:0] PEManager_15U_GetWeightAddr_else_acc_3_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
  reg [63:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
  reg [63:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
  reg [63:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
  reg [17:0] Datapath_for_3_ProductSum_for_acc_3_1;
  reg [15:0] act_port_reg_data_239_224_sva_dfm_1_1;
  reg [15:0] act_port_reg_data_207_192_sva_dfm_1_1;
  reg [15:0] act_port_reg_data_175_160_sva_dfm_1_1;
  reg [15:0] act_port_reg_data_143_128_sva_dfm_1_1;
  reg [15:0] act_port_reg_data_111_96_sva_dfm_1_1;
  reg [15:0] act_port_reg_data_47_32_sva_dfm_1_1;
  reg [15:0] act_port_reg_data_15_0_sva_dfm_1_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  reg [14:0] pe_manager_base_weight_sva_dfm_3_1;
  reg [14:0] pe_manager_base_input_sva_dfm_3_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_55_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1;
  reg [7:0] weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1;
  reg [7:0] weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_2;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1;
  reg weight_mem_run_3_for_5_and_162_itm_1;
  reg weight_mem_run_3_for_5_and_163_itm_1;
  reg weight_mem_run_3_for_5_and_164_itm_1;
  reg weight_mem_run_3_for_5_and_164_itm_2;
  reg weight_mem_run_3_for_5_and_165_itm_1;
  reg weight_mem_run_3_for_5_and_166_itm_1;
  reg weight_mem_run_3_for_5_and_167_itm_1;
  reg weight_mem_run_3_for_5_and_168_itm_1;
  reg weight_mem_run_3_for_5_and_8_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
  reg weight_mem_run_3_for_5_and_20_itm_1;
  reg weight_mem_run_3_for_5_and_20_itm_2;
  reg weight_mem_run_3_for_5_and_22_itm_1;
  reg weight_mem_run_3_for_5_and_23_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1;
  reg weight_mem_run_3_for_5_and_28_itm_1;
  reg weight_mem_run_3_for_5_and_30_itm_1;
  reg weight_mem_run_3_for_5_and_30_itm_2;
  reg weight_mem_run_3_for_5_and_31_itm_1;
  reg weight_mem_run_3_for_5_and_31_itm_2;
  reg weight_mem_run_3_for_5_and_79_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1;
  reg weight_mem_run_3_for_5_and_84_itm_1;
  reg weight_mem_run_3_for_5_and_86_itm_1;
  reg weight_mem_run_3_for_5_and_86_itm_2;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2;
  reg weight_mem_run_3_for_5_and_92_itm_1;
  reg weight_mem_run_3_for_5_and_92_itm_2;
  reg weight_mem_run_3_for_5_and_94_itm_1;
  reg weight_mem_run_3_for_5_and_95_itm_1;
  reg weight_mem_run_3_for_5_and_95_itm_2;
  reg weight_mem_run_3_for_5_and_96_itm_1;
  reg weight_mem_run_3_for_5_and_103_itm_1;
  reg weight_mem_run_3_for_5_and_103_itm_2;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2;
  reg weight_mem_run_3_for_5_and_144_itm_1;
  reg weight_mem_run_3_for_5_and_150_itm_1;
  reg weight_mem_run_3_for_5_and_150_itm_2;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1;
  reg weight_mem_run_3_for_5_and_156_itm_1;
  reg weight_mem_run_3_for_5_and_156_itm_2;
  reg weight_mem_run_3_for_5_and_158_itm_1;
  reg weight_mem_run_3_for_5_and_159_itm_1;
  reg [18:0] ProductSum_for_acc_22_itm_1;
  wire [19:0] nl_ProductSum_for_acc_22_itm_1;
  reg [14:0] PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1;
  reg while_if_mux_19_itm_1;
  reg PECore_PushAxiRsp_mux_10_itm_1;
  reg PECore_PushAxiRsp_mux_13_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
  reg [55:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_1_63_8;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0;
  reg [31:0] input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0;
  reg [31:0] input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_3_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0;
  wire PECore_PushAxiRsp_if_else_mux_13_mx0w2;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_39_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_38_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_37_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0;
  wire weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_2_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0;
  wire [14:0] weight_read_addrs_1_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_3_lpi_1_dfm_1_1;
  wire [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_5_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_7_lpi_1_dfm_1_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  wire [7:0] pe_config_output_counter_sva_mx1;
  wire pe_config_is_zero_first_sva_mx1;
  wire pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  wire [15:0] act_port_reg_data_79_64_sva_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
  wire [15:0] act_port_reg_data_15_0_sva_mx1;
  wire [15:0] act_port_reg_data_47_32_sva_mx1;
  wire [15:0] act_port_reg_data_111_96_sva_mx1;
  wire [15:0] act_port_reg_data_143_128_sva_mx1;
  wire [15:0] act_port_reg_data_175_160_sva_mx1;
  wire [15:0] act_port_reg_data_207_192_sva_mx1;
  wire [15:0] act_port_reg_data_239_224_sva_mx1;
  wire [63:0] input_mem_banks_bank_a_0_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_1_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_2_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_3_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_4_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_5_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_6_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_7_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_8_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_9_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_10_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_11_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_12_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_13_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_14_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_15_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_16_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_17_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_18_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_19_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_20_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_21_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_22_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_23_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_24_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_25_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_26_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_27_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_28_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_29_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_30_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_31_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_32_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_33_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_34_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_35_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_36_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_37_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_38_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_39_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_40_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_41_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_42_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_43_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_44_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_45_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_46_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_47_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_48_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_49_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_50_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_51_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_52_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_53_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_54_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_55_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_56_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_57_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_58_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_59_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_60_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_61_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_62_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_63_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_64_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_65_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_66_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_67_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_68_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_69_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_70_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_71_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_72_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_73_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_74_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_75_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_76_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_77_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_78_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_79_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_80_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_81_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_82_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_83_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_84_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_85_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_86_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_87_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_88_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_89_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_90_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_91_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_92_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_93_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_94_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_95_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_96_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_97_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_98_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_99_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_100_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_101_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_102_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_103_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_104_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_105_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_106_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_107_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_108_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_109_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_110_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_111_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_112_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_113_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_114_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_115_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_116_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_117_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_118_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_119_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_120_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_121_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_122_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_123_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_124_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_125_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_126_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_127_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_128_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_129_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_130_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_131_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_132_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_133_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_134_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_135_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_136_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_137_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_138_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_139_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_140_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_141_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_142_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_143_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_144_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_145_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_146_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_147_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_148_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_149_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_150_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_151_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_152_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_153_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_154_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_155_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_156_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_157_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_158_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_159_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_160_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_161_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_162_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_163_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_164_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_165_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_166_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_167_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_168_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_169_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_170_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_171_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_172_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_173_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_174_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_175_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_176_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_177_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_178_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_179_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_180_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_181_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_182_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_183_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_184_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_185_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_186_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_187_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_188_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_189_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_190_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_191_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_192_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_193_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_194_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_195_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_196_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_197_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_198_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_199_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_200_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_201_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_202_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_203_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_204_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_205_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_206_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_207_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_208_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_209_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_210_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_211_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_212_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_213_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_214_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_215_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_216_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_217_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_218_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_219_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_220_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_221_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_222_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_223_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_224_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_225_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_226_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_227_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_228_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_229_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_230_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_231_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_232_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_233_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_234_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_235_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_236_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_237_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_238_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_239_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_240_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_241_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_242_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_243_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_244_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_245_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_246_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_247_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_248_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_249_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_250_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_251_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_252_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_253_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_254_sva_dfm_2_mx0w0;
  wire [63:0] input_mem_banks_bank_a_255_sva_dfm_2_mx0w0;
  wire PECore_PushAxiRsp_if_else_mux_10_mx0w2;
  wire [6:0] rva_out_reg_data_62_56_sva_dfm_6_mx1;
  wire [3:0] rva_out_reg_data_35_32_sva_dfm_6_mx1;
  wire PECore_PushAxiRsp_mux_13_itm_1_mx0c1;
  wire [14:0] pe_manager_base_input_sva_mx2;
  wire PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  wire [7:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1;
  wire weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_4;
  wire while_and_1129_cse_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14;
  wire rva_out_reg_data_63_sva_dfm_7;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_257_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_255_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_256_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_254_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_255_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_253_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_254_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_252_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_253_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_251_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_252_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_250_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_251_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_249_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_250_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_248_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_249_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_247_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_248_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_246_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_247_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_245_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_246_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_244_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_245_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_243_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_244_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_242_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_243_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_241_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_242_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_240_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_241_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_239_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_240_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_238_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_239_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_237_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_238_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_236_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_237_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_235_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_236_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_234_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_235_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_233_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_234_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_232_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_233_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_231_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_232_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_230_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_231_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_229_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_230_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_228_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_229_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_227_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_228_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_226_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_227_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_225_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_226_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_224_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_225_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_223_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_224_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_222_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_223_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_221_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_222_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_220_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_221_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_219_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_220_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_218_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_219_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_217_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_218_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_216_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_217_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_215_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_216_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_214_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_215_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_213_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_214_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_212_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_213_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_211_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_212_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_210_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_211_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_209_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_210_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_208_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_209_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_207_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_208_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_206_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_207_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_205_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_206_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_204_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_205_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_203_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_204_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_202_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_203_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_201_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_202_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_200_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_201_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_199_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_200_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_198_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_199_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_197_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_198_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_196_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_197_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_195_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_196_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_194_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_195_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_193_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_194_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_192_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_193_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_191_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_192_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_190_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_191_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_189_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_190_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_188_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_189_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_187_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_188_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_186_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_187_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_185_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_186_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_184_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_185_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_183_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_184_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_182_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_183_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_181_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_182_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_180_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_181_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_179_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_180_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_178_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_179_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_177_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_178_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_176_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_177_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_175_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_176_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_174_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_175_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_173_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_174_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_172_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_173_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_171_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_172_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_170_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_171_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_169_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_170_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_168_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_169_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_167_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_168_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_166_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_167_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_165_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_166_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_164_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_165_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_163_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_164_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_162_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_163_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_161_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_162_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_160_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_161_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_159_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_160_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_158_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_159_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_157_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_158_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_156_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_157_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_155_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_156_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_154_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_155_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_153_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_154_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_152_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_153_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_151_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_152_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_150_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_151_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_149_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_150_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_148_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_149_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_147_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_148_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_146_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_147_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_145_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_146_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_144_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_145_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_143_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_144_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_142_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_143_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_141_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_142_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_140_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_141_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_139_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_140_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_138_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_139_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_137_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_138_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_136_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_137_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_135_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_136_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_134_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_135_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_133_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_134_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_132_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_133_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_131_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_132_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_130_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_131_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_129_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_130_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_128_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_129_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_127_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_128_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_126_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_127_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_125_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_126_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_124_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_125_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_123_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_124_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_122_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_123_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_121_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_122_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_120_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_121_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_119_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_120_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_118_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_119_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_117_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_118_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_116_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_117_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_115_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_116_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_114_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_115_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_113_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_114_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_112_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_113_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_111_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_112_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_110_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_111_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_109_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_110_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_108_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_109_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_107_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_108_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_106_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_107_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_105_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_106_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_104_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_105_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_103_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_104_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_102_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_103_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_101_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_102_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_100_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_101_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_99_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_100_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_98_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_99_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_97_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_98_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_96_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_97_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_95_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_96_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_94_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_95_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_93_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_94_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_92_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_93_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_91_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_92_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_90_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_91_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_89_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_90_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_88_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_89_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_87_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_88_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_86_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_87_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_85_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_86_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_84_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_85_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_83_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_84_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_82_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_83_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_81_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_82_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_80_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_81_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_79_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_80_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_78_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_79_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_77_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_78_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_76_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_77_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_75_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_76_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_74_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_75_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_73_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_74_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_72_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_73_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_71_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_72_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_70_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_71_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_69_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_70_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_68_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_69_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_67_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_68_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_66_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_67_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_65_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_66_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_64_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_65_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_63_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_64_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_62_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_63_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_61_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_62_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_60_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_61_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_59_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_60_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_58_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_59_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_57_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_58_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_56_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_57_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_55_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_56_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_54_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_55_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_53_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_54_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_52_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_53_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_51_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_52_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_50_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_51_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_49_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_50_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_48_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_49_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_47_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_48_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_46_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_47_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_45_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_46_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_44_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_45_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_43_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_44_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_42_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_43_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_41_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_42_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_40_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_41_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_39_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_40_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_38_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_39_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_37_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_38_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_36_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_37_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_35_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_36_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_34_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_35_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_33_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_34_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_32_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_33_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_31_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_32_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_30_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_31_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_29_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_30_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_28_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_29_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_27_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_28_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_26_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_27_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_25_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_26_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_24_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_25_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_23_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_24_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_22_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_23_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_21_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_22_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_20_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_21_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_19_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_20_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_18_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_19_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_17_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_18_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_16_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_17_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_15_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_16_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_14_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_15_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_13_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_14_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_12_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_13_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_11_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_12_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_10_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_11_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_9_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_10_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_8_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_9_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_7_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_8_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_6_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_7_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_5_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_6_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_4_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_5_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_3_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_4_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_2_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_3_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_1_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_2_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_tmp_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
  wire PECore_PushAxiRsp_if_asn_55;
  wire PECore_PushAxiRsp_if_asn_57;
  wire PECore_PushAxiRsp_if_asn_59;
  wire weight_mem_run_3_for_5_asn_308;
  wire weight_mem_run_3_for_5_asn_310;
  wire weight_mem_run_3_for_5_asn_312;
  wire weight_mem_run_3_for_5_asn_314;
  wire weight_mem_run_3_for_5_asn_316;
  wire weight_mem_run_3_for_5_asn_318;
  wire weight_mem_run_3_for_5_asn_320;
  wire weight_mem_run_3_for_5_asn_322;
  wire weight_mem_run_3_for_5_asn_324;
  wire weight_mem_run_3_for_5_asn_326;
  wire weight_mem_run_3_for_5_asn_328;
  wire weight_mem_run_3_for_5_asn_330;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56;
  wire PECore_PushAxiRsp_if_asn_61;
  wire PECore_PushAxiRsp_if_asn_63;
  wire PECore_PushAxiRsp_if_asn_65;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98;
  wire weight_mem_run_3_for_5_and_166;
  wire weight_mem_run_3_for_5_and_168;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100;
  wire weight_mem_run_3_for_5_and_172;
  wire weight_mem_run_3_for_5_and_174;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54;
  wire [7:0] pe_manager_base_input_sva_mx1_7_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0;
  wire PECore_PushAxiRsp_if_mux1h_15;
  wire PECore_PushAxiRsp_if_mux1h_17;
  wire [7:0] weight_port_read_out_data_3_4_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_3_5_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_5_6_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_5_7_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_5_4_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_5_5_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_5_2_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_5_3_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_5_0_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_5_1_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_3_6_sva_dfm_3;
  wire [7:0] weight_port_read_out_data_3_7_sva_dfm_3;
  reg reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_162_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_163_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_165_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_166_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_167_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_168_itm_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse;
  reg reg_rva_in_reg_rw_sva_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse;
  wire weight_mem_run_3_for_5_and_222_ssc;
  reg weight_mem_run_3_for_5_mux_17_itm_1_7;
  wire weight_port_read_out_data_and_94_ssc;
  reg weight_port_read_out_data_0_3_sva_dfm_1_7;
  wire weight_mem_banks_load_store_for_else_and_1_ssc;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7_4;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0;
  wire weight_mem_banks_load_store_for_else_and_17_ssc;
  reg [1:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6;
  reg [5:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0;
  wire weight_mem_banks_load_store_for_else_and_7_ssc;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0;
  reg weight_port_read_out_data_0_3_sva_dfm_2_7;
  reg weight_port_read_out_data_0_2_sva_dfm_2_7;
  wire weight_port_read_out_data_0_1_sva_dfm_mx0w1_7;
  wire [6:0] weight_port_read_out_data_0_1_sva_dfm_mx0w1_6_0;
  wire and_936_ssc;
  wire weight_port_read_out_data_0_0_sva_dfm_mx0w1_7;
  wire [6:0] weight_port_read_out_data_0_0_sva_dfm_mx0w1_6_0;
  wire and_945_ssc;
  wire weight_port_read_out_data_0_2_sva_dfm_mx0w2_7;
  wire weight_port_read_out_data_0_2_sva_dfm_mx0w2_6;
  wire [5:0] weight_port_read_out_data_0_2_sva_dfm_mx0w2_5_0;
  wire weight_port_read_out_data_0_3_sva_dfm_mx0w0_7;
  wire [2:0] weight_port_read_out_data_0_3_sva_dfm_mx0w0_6_4;
  wire [3:0] weight_port_read_out_data_0_3_sva_dfm_mx0w0_3_0;
  wire [3:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_7_4;
  wire [3:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_3_0;
  wire weight_port_read_out_data_0_7_sva_dfm_3_7;
  wire [6:0] weight_port_read_out_data_0_7_sva_dfm_3_6_0;
  wire and_972_ssc;
  wire and_973_ssc;
  wire and_974_ssc;
  wire and_975_ssc;
  wire and_976_ssc;
  wire and_977_ssc;
  wire and_978_ssc;
  wire nor_431_ssc;
  wire [3:0] weight_port_read_out_data_0_5_sva_dfm_3_7_4;
  wire [3:0] weight_port_read_out_data_0_5_sva_dfm_3_3_0;
  wire and_981_ssc;
  wire and_984_ssc;
  wire and_985_ssc;
  wire weight_port_read_out_data_0_4_sva_dfm_3_7;
  wire weight_port_read_out_data_0_4_sva_dfm_3_6;
  wire [5:0] weight_port_read_out_data_0_4_sva_dfm_3_5_0;
  reg weight_port_read_out_data_0_2_sva_dfm_3_rsp_0;
  reg weight_port_read_out_data_0_3_sva_dfm_3_rsp_0;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd;
  reg weight_port_read_out_data_0_1_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_1_sva_dfm_2_6_0;
  reg weight_port_read_out_data_0_3_sva_dfm_2_7_1;
  reg [2:0] weight_port_read_out_data_0_3_sva_dfm_2_6_4;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_2_3_0;
  reg weight_port_read_out_data_0_2_sva_dfm_2_7_1;
  reg weight_port_read_out_data_0_2_sva_dfm_2_6;
  reg [5:0] weight_port_read_out_data_0_2_sva_dfm_2_5_0;
  reg [3:0] weight_port_read_out_data_0_5_sva_dfm_2_7_4;
  reg [3:0] weight_port_read_out_data_0_5_sva_dfm_2_3_0;
  reg weight_port_read_out_data_0_4_sva_dfm_2_7;
  reg weight_port_read_out_data_0_4_sva_dfm_2_6;
  reg [5:0] weight_port_read_out_data_0_4_sva_dfm_2_5_0;
  reg weight_port_read_out_data_0_7_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_7_sva_dfm_2_6_0;
  wire weight_port_read_out_data_and_1_ssc;
  reg [3:0] weight_port_read_out_data_0_6_sva_dfm_2_7_4;
  reg [3:0] weight_port_read_out_data_0_6_sva_dfm_2_3_0;
  reg input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_7;
  reg [6:0] input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_6_0;
  wire input_mem_banks_read_1_read_data_and_ssc;
  reg input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_7;
  reg [6:0] input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_6_0;
  reg weight_port_read_out_data_0_0_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_0_sva_dfm_2_6_0;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_1_7_4;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_1_3_0;
  reg [2:0] rva_out_reg_data_46_40_sva_dfm_4_1_6_4;
  reg [3:0] rva_out_reg_data_46_40_sva_dfm_4_1_3_0;
  reg rva_out_reg_data_39_36_sva_dfm_4_1_3;
  reg rva_out_reg_data_39_36_sva_dfm_4_1_2;
  reg [1:0] rva_out_reg_data_39_36_sva_dfm_4_1_1_0;
  reg weight_mem_run_3_for_5_mux_17_itm_1_6;
  reg [5:0] weight_mem_run_3_for_5_mux_17_itm_1_5_0;
  reg [2:0] weight_port_read_out_data_0_3_sva_dfm_1_6_4;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_1_3_0;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_5_a_mx1_7;
  wire [6:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_a_mx1_6_0;
  wire weight_port_read_out_data_0_0_sva_dfm_3_7;
  wire [6:0] weight_port_read_out_data_0_0_sva_dfm_3_6_0;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_7;
  wire [2:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_6_4;
  wire [3:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_3_0;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_7;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_6;
  wire [5:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_5_0;
  wire weight_mem_run_3_for_5_and_190_ssc;
  wire weight_mem_run_3_for_5_and_191_ssc;
  wire weight_mem_run_3_for_5_and_192_ssc;
  wire weight_mem_run_3_for_5_and_193_ssc;
  wire weight_mem_run_3_for_5_and_194_ssc;
  wire weight_mem_run_3_for_5_and_195_ssc;
  wire [3:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_a_mx1_7_4;
  wire [3:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_a_mx1_3_0;
  wire weight_mem_run_3_for_5_and_187_ssc;
  wire weight_mem_run_3_for_5_and_188_ssc;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_7;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_6;
  wire [5:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_5_0;
  wire weight_mem_run_3_for_5_and_ssc;
  wire weight_mem_run_3_for_5_and_179_ssc;
  wire weight_mem_run_3_for_5_and_180_ssc;
  wire weight_mem_run_3_for_5_and_181_ssc;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_8_a_mx1_7;
  wire [6:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_a_mx1_6_0;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_2_7_4;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_2_3_0;
  reg [2:0] rva_out_reg_data_46_40_sva_dfm_4_2_6_4;
  reg [3:0] rva_out_reg_data_46_40_sva_dfm_4_2_3_0;
  reg rva_out_reg_data_39_36_sva_dfm_4_2_3;
  reg rva_out_reg_data_39_36_sva_dfm_4_2_2;
  reg [1:0] rva_out_reg_data_39_36_sva_dfm_4_2_1_0;
  reg weight_port_read_out_data_0_3_sva_dfm_5_7;
  reg weight_port_read_out_data_0_1_sva_dfm_2_7_1;
  reg [6:0] weight_port_read_out_data_0_1_sva_dfm_2_6_0_1;
  wire weight_port_read_out_data_and_90_ssc;
  reg weight_port_read_out_data_0_0_sva_dfm_2_7_1;
  reg [6:0] weight_port_read_out_data_0_0_sva_dfm_2_6_0_1;
  reg rva_out_reg_data_15_9_sva_dfm_7_6;
  reg [5:0] rva_out_reg_data_15_9_sva_dfm_7_5_0;
  reg [2:0] rva_out_reg_data_23_17_sva_dfm_5_6_4;
  reg [3:0] rva_out_reg_data_23_17_sva_dfm_5_3_0;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_6;
  wire [3:0] rva_out_reg_data_55_48_sva_dfm_6_mx1_7_4;
  wire [3:0] rva_out_reg_data_55_48_sva_dfm_6_mx1_3_0;
  wire [2:0] rva_out_reg_data_46_40_sva_dfm_6_mx1_6_4;
  wire [3:0] rva_out_reg_data_46_40_sva_dfm_6_mx1_3_0;
  wire rva_out_reg_data_39_36_sva_dfm_6_mx1_3;
  wire rva_out_reg_data_39_36_sva_dfm_6_mx1_2;
  wire [1:0] rva_out_reg_data_39_36_sva_dfm_6_mx1_1_0;
  reg [2:0] weight_port_read_out_data_0_3_sva_dfm_2_6_4_1;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_2_3_0_1;
  reg weight_port_read_out_data_0_2_sva_dfm_2_6_1;
  reg [5:0] weight_port_read_out_data_0_2_sva_dfm_2_5_0_1;
  wire rva_out_reg_data_and_14_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_2_cse;
  wire rva_out_reg_data_and_17_cse;
  wire input_mem_banks_read_read_data_and_cse;
  wire weight_port_read_out_data_and_64_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_cse;
  wire act_port_reg_data_and_cse;
  wire rva_in_reg_rw_and_cse;
  wire weight_mem_run_3_for_aelse_and_cse;
  wire weight_mem_banks_read_1_read_data_and_8_cse;
  wire weight_mem_run_3_for_aelse_and_1_cse;
  wire weight_port_read_out_data_and_71_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_101_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_113_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_49_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_55_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_61_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_67_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_73_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_79_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_85_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_91_cse;
  wire weight_read_addrs_and_9_cse;
  wire weight_write_data_data_and_cse;
  wire weight_mem_write_arbxbar_xbar_for_1_for_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse;
  wire PECore_RunFSM_switch_lp_and_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_15_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_22_cse;
  wire Arbiter_8U_Roundrobin_pick_and_75_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_23_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_64_cse;
  wire weight_write_data_data_and_8_cse;
  wire rva_in_reg_rw_and_6_cse;
  wire PECore_UpdateFSM_switch_lp_and_9_cse;
  wire state_and_cse;
  wire PECore_PushOutput_if_and_cse;
  wire PECore_RunMac_if_and_cse;
  wire weight_mem_banks_load_store_for_else_and_cse;
  wire weight_mem_banks_load_store_for_else_and_6_cse;
  wire weight_mem_banks_load_store_for_else_and_10_cse;
  wire weight_mem_banks_load_store_for_else_and_14_cse;
  wire weight_mem_banks_load_store_for_else_and_9_cse;
  wire weight_mem_banks_load_store_for_else_and_19_cse;
  wire weight_mem_banks_load_store_for_else_and_16_cse;
  wire weight_read_addrs_and_19_cse;
  wire while_if_and_11_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_24_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_122_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_74_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_79_cse;
  wire weight_port_read_out_data_and_79_cse;
  wire input_mem_banks_read_read_data_and_9_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse;
  wire while_if_and_15_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_7_cse;
  wire while_if_and_6_cse;
  wire rva_out_reg_data_and_24_cse;
  wire input_read_req_valid_and_1_cse;
  wire ProductSum_for_and_cse;
  wire weight_port_read_out_data_and_86_cse;
  wire rva_in_reg_rw_and_7_cse;
  wire PECore_RunMac_if_and_1_cse;
  wire input_mem_banks_read_read_data_and_18_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_11_cse;
  wire while_if_and_7_cse;
  wire rva_out_reg_data_and_34_cse;
  wire input_read_req_valid_and_2_cse;
  wire PECore_RunScale_if_and_1_cse;
  wire PECore_RunMac_if_and_2_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_15_cse;
  wire while_if_and_8_cse;
  wire rva_out_reg_data_and_42_cse;
  wire input_read_req_valid_and_3_cse;
  wire PECore_RunMac_if_and_3_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse;
  wire PECore_RunScale_if_and_2_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_19_cse;
  wire rva_out_reg_data_and_51_cse;
  wire input_read_req_valid_and_4_cse;
  wire rva_out_reg_data_and_56_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse;
  wire PECore_RunScale_if_and_3_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_23_cse;
  wire PECore_RunMac_if_and_6_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_23_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_27_cse;
  wire rva_out_reg_data_and_62_cse;
  wire rva_out_reg_data_and_65_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_28_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_31_cse;
  wire rva_out_reg_data_and_70_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_33_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_35_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse;
  wire while_if_and_16_cse;
  wire rva_out_reg_data_and_85_cse;
  wire rva_out_reg_data_and_61_cse;
  reg weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
  reg [6:0] weight_port_read_out_data_0_0_sva_dfm_3_rsp_1;
  reg weight_port_read_out_data_0_1_sva_dfm_3_rsp_0;
  reg [6:0] weight_port_read_out_data_0_1_sva_dfm_3_rsp_1;
  reg [2:0] rva_out_reg_data_23_17_sva_dfm_6_rsp_0;
  reg [3:0] rva_out_reg_data_23_17_sva_dfm_6_rsp_1;
  reg rva_out_reg_data_15_9_sva_dfm_8_rsp_0;
  reg [5:0] rva_out_reg_data_15_9_sva_dfm_8_rsp_1;
  reg rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0;
  reg rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1;
  reg [1:0] rva_out_reg_data_39_36_sva_dfm_4_3_rsp_2;
  reg [2:0] rva_out_reg_data_46_40_sva_dfm_4_3_rsp_0;
  reg [3:0] rva_out_reg_data_46_40_sva_dfm_4_3_rsp_1;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_3_rsp_0;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_3_rsp_1;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_6_rsp_0;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_6_rsp_1;
  reg [2:0] rva_out_reg_data_46_40_sva_dfm_6_rsp_0;
  reg [3:0] rva_out_reg_data_46_40_sva_dfm_6_rsp_1;
  reg rva_out_reg_data_39_36_sva_dfm_6_rsp_0;
  reg rva_out_reg_data_39_36_sva_dfm_6_rsp_1;
  reg [1:0] rva_out_reg_data_39_36_sva_dfm_6_rsp_2;
  reg weight_port_read_out_data_0_2_sva_dfm_3_rsp_1_rsp_0;
  reg [5:0] weight_port_read_out_data_0_2_sva_dfm_3_rsp_1_rsp_1;
  reg [2:0] weight_port_read_out_data_0_3_sva_dfm_3_rsp_1_rsp_0;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_3_rsp_1_rsp_1;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd;
  reg [5:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd;
  reg [5:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_1_ftd;
  reg [4:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_1_ftd_1;
  reg [2:0] reg_rva_out_reg_data_23_17_sva_dfm_7_ftd;
  reg [3:0] reg_rva_out_reg_data_23_17_sva_dfm_7_ftd_1;
  reg reg_rva_out_reg_data_15_9_sva_dfm_9_ftd;
  reg [5:0] reg_rva_out_reg_data_15_9_sva_dfm_9_ftd_1;
  reg [2:0] reg_weight_port_read_out_data_0_3_sva_dfm_4_1_ftd;
  reg [3:0] reg_weight_port_read_out_data_0_3_sva_dfm_4_1_ftd_1;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1;
  reg [1:0] reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_2;
  reg [2:0] reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd;
  reg [3:0] reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd_1;
  reg [3:0] reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd;
  reg [3:0] reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd_1;
  wire PECore_PushAxiRsp_if_mux1h_14_6;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_5_7_4;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_5_3_0;
  reg [2:0] rva_out_reg_data_46_40_sva_dfm_4_5_6_4;
  reg [3:0] rva_out_reg_data_46_40_sva_dfm_4_5_3_0;
  reg rva_out_reg_data_39_36_sva_dfm_4_5_3;
  reg rva_out_reg_data_39_36_sva_dfm_4_5_2;
  reg [1:0] rva_out_reg_data_39_36_sva_dfm_4_5_1_0;
  reg rva_out_reg_data_23_17_sva_dfm_6_6;
  reg rva_out_reg_data_15_9_sva_dfm_10_6;
  reg [5:0] rva_out_reg_data_15_9_sva_dfm_10_5_0;
  reg [2:0] rva_out_reg_data_23_17_sva_dfm_8_6_4;
  reg [3:0] rva_out_reg_data_23_17_sva_dfm_8_3_0;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_6;
  reg [5:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_5_0;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_6;
  reg [5:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_5_0;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_5_0_rsp_0;
  reg [4:0] weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_5_0_rsp_1;
  reg [2:0] weight_port_read_out_data_0_3_sva_dfm_5_6_0_rsp_0;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_5_6_0_rsp_1;
  wire PECore_PushAxiRsp_if_mux1h_10_6;
  wire [5:0] PECore_PushAxiRsp_if_mux1h_10_5_0;
  wire PECore_PushAxiRsp_if_mux1h_12_6;
  wire [5:0] PECore_PushAxiRsp_if_mux1h_12_5_0;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_16_5_3;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_16_2_0;
  wire PECore_PushAxiRsp_if_mux1h_14_5;
  wire PECore_PushAxiRsp_if_mux1h_14_4;
  wire [3:0] PECore_PushAxiRsp_if_mux1h_14_3_0;
  reg [2:0] rva_out_reg_data_30_25_sva_dfm_6_5_3;
  reg [2:0] rva_out_reg_data_30_25_sva_dfm_6_2_0;
  reg rva_out_reg_data_15_9_sva_dfm_6_6;
  reg [5:0] rva_out_reg_data_15_9_sva_dfm_6_5_0;
  reg rva_out_reg_data_7_1_sva_dfm_6_6;
  reg [5:0] rva_out_reg_data_7_1_sva_dfm_6_5_0;
  reg rva_out_reg_data_23_17_sva_dfm_6_5;
  reg rva_out_reg_data_23_17_sva_dfm_6_4;
  reg [3:0] rva_out_reg_data_23_17_sva_dfm_6_3_0;
  wire or_dcpl_308;
  wire or_dcpl_312;
  wire or_dcpl_330;
  wire and_dcpl_719;
  wire or_dcpl_345;
  wire or_dcpl_350;
  wire or_dcpl_355;
  wire or_dcpl_382;
  wire and_dcpl_811;
  wire [7:0] PEManager_15U_GetInputAddr_acc_tmp;
  wire [8:0] nl_PEManager_15U_GetInputAddr_acc_tmp;
  wire or_tmp_1863;
  wire and_1010_cse;
  wire and_1019_cse;
  wire mux_340_cse;
  wire and_1043_cse;
  wire xor_7_cse;
  wire and_1083_cse;
  wire xor_13_cse;
  wire or_835_cse;
  wire or_228_cse_1;
  wire and_1169_cse;
  wire and_1197_cse;
  wire and_1231_cse;
  wire and_1258_cse;
  wire or_898_cse;
  wire nand_247_cse;
  wire nand_248_cse;
  wire nand_250_cse;
  wire nand_254_cse;
  wire nand_262_cse;
  wire and_1792_cse;
  wire mux_85_cse;
  wire nor_718_cse;
  wire and_1109_cse;
  wire and_1884_cse;
  wire nor_690_cse;
  wire nor_695_cse;
  wire and_2190_cse;
  wire and_1018_cse;
  wire and_1030_cse;
  wire and_1054_cse;
  wire and_1059_cse;
  wire and_1044_cse;
  wire mux_365_cse;
  wire mux_387_cse;
  wire mux_389_cse;
  wire mux_403_cse;
  wire mux_415_cse;
  wire mux_417_cse;
  wire and_1801_cse;
  wire and_1831_cse;
  wire and_1840_cse;
  wire and_1835_cse;
  wire or_2320_cse;
  reg reg_rva_out_reg_data_30_25_sva_dfm_7_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  reg reg_act_port_reg_data_15_0_sva_dfm_1_1_enexo;
  reg reg_act_port_reg_data_239_224_sva_dfm_1_1_enexo;
  reg reg_act_port_reg_data_47_32_sva_dfm_1_1_enexo;
  reg reg_act_port_reg_data_207_192_sva_dfm_1_1_enexo;
  reg reg_act_port_reg_data_175_160_sva_dfm_1_1_enexo;
  reg reg_act_port_reg_data_111_96_sva_dfm_1_1_enexo;
  reg reg_act_port_reg_data_143_128_sva_dfm_1_1_enexo;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_000000;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo;
  reg reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo_1;
  reg reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2;
  reg reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_manager_base_input_enexo;
  reg reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_config_num_output_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  reg reg_rva_in_reg_data_sva_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_3_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_6_1_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_8_1_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_3_2_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_3_1_enexo;
  reg reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_1;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_2;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_3;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0_enexo;
  reg reg_input_mem_banks_bank_a_189_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_208_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_21_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_188_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_22_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_249_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_221_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_113_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_88_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_13_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_27_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_72_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_46_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_132_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_155_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_157_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_243_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_149_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_49_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_220_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_90_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_83_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_81_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_241_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_50_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_96_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_123_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_12_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_250_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_248_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_246_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_95_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_255_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_17_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_235_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_214_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_251_sva_dfm_2_enexo;
  reg reg_input_read_addrs_sva_1_1_enexo;
  reg reg_input_mem_banks_bank_a_231_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_104_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_142_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_109_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_36_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_8_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_19_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_181_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_177_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_191_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_4_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_204_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_53_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_116_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_139_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_110_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_136_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_91_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_55_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_68_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_224_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_223_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_93_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_75_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_135_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_150_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_108_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_169_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_52_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_240_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_213_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_121_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_14_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_192_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_194_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_172_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_117_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_197_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_71_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_31_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_41_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_158_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_58_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_76_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_24_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_65_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_40_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_30_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_151_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_44_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_107_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_1_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_39_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_61_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_137_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_222_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_165_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_94_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_254_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_207_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_47_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_89_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_228_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_234_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_193_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_187_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_45_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_112_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_11_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_66_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_15_sva_dfm_2_enexo;
  reg reg_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1_enexo;
  reg reg_input_mem_banks_bank_a_184_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_103_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_124_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_182_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_247_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_84_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_167_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_148_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_227_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_232_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_186_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_253_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_105_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_101_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_7_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_5_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_201_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_236_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_195_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_62_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_92_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_18_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_35_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_210_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_106_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_70_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_126_sva_dfm_2_enexo;
  reg reg_input_mem_banks_read_read_data_sva_1_enexo;
  reg reg_input_mem_banks_bank_a_3_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_97_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_252_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_77_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_57_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_217_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_163_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_16_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_42_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_219_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_225_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_120_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_63_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_229_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_176_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_54_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_74_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_80_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_78_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_140_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_153_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_174_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_156_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_202_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_238_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_67_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_87_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_147_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_170_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_2_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_29_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_183_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_166_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_33_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_134_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_162_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_159_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_51_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_152_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_173_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_179_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_180_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_144_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_209_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_48_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_160_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_203_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_20_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_43_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_237_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_102_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_111_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_129_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_100_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_10_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_145_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_239_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_196_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_56_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_154_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_141_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_245_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_128_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_164_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_175_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_69_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_6_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_125_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_127_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_82_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_25_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_226_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_138_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_133_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_37_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_242_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_171_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_216_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_206_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_9_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_32_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_86_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_122_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_26_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_190_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_199_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_73_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_79_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_114_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_131_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_198_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_98_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_168_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_146_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_211_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_233_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_115_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_215_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_212_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_200_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_143_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_185_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_23_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_205_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_99_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_38_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_230_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_218_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_244_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_161_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_60_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_130_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_178_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_119_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_118_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_34_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_28_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_85_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_64_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_59_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_0_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_4_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_1_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_1_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_5_1_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_7_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_2_1_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo;
  reg reg_weight_mem_run_3_for_5_mux_17_itm_1_2_enexo;
  reg reg_input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_1_enexo;
  reg reg_input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_1_1_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_2_2_enexo;
  reg reg_weight_mem_run_3_for_5_mux_17_itm_1_2_enexo_1;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo_1;
  reg reg_rva_out_reg_data_15_9_sva_dfm_9_1_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_7_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_4_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_4_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_4_1_enexo;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_1_enexo;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_1_enexo;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_2_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_4_2_enexo;
  wire rva_out_reg_data_and_90_enex5;
  wire rva_out_reg_data_and_91_enex5;
  wire rva_out_reg_data_and_92_enex5;
  wire input_mem_banks_read_read_data_and_31_enex5;
  wire input_mem_banks_read_read_data_and_32_enex5;
  wire input_mem_banks_read_read_data_and_33_enex5;
  wire input_mem_banks_read_read_data_and_34_enex5;
  wire act_port_reg_data_and_30_enex5;
  wire act_port_reg_data_and_31_enex5;
  wire act_port_reg_data_and_32_enex5;
  wire act_port_reg_data_and_33_enex5;
  wire act_port_reg_data_and_34_enex5;
  wire act_port_reg_data_and_35_enex5;
  wire act_port_reg_data_and_36_enex5;
  wire weight_port_read_out_data_and_enex5;
  wire input_mem_banks_read_1_read_data_and_2_enex5;
  wire weight_read_addrs_and_7_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5;
  wire weight_write_data_data_and_24_enex5;
  wire weight_write_data_data_and_25_enex5;
  wire weight_write_data_data_and_26_enex5;
  wire weight_write_data_data_and_27_enex5;
  wire weight_write_data_data_and_28_enex5;
  wire weight_write_data_data_and_29_enex5;
  wire weight_write_data_data_and_30_enex5;
  wire weight_write_data_data_and_31_enex5;
  wire weight_write_addrs_and_enex5;
  wire weight_write_data_data_and_32_enex5;
  wire weight_write_data_data_and_33_enex5;
  wire weight_write_data_data_and_34_enex5;
  wire weight_write_data_data_and_35_enex5;
  wire weight_write_data_data_and_36_enex5;
  wire weight_write_data_data_and_37_enex5;
  wire weight_write_data_data_and_38_enex5;
  wire weight_write_data_data_and_39_enex5;
  wire weight_write_addrs_and_2_enex5;
  wire weight_read_addrs_and_28_enex5;
  wire pe_config_UpdateManagerCounter_if_if_and_enex5;
  wire weight_read_addrs_and_29_enex5;
  wire PEManager_15U_PEManagerWrite_and_enex5;
  wire weight_port_read_out_data_and_95_enex5;
  wire input_mem_banks_read_read_data_and_35_enex5;
  wire weight_port_read_out_data_and_96_enex5;
  wire input_mem_banks_read_read_data_and_36_enex5;
  wire weight_port_read_out_data_and_97_enex5;
  wire input_mem_banks_read_read_data_and_37_enex5;
  wire input_mem_banks_read_read_data_and_38_enex5;
  wire input_mem_banks_read_1_read_data_and_3_enex5;
  wire rva_out_reg_data_and_93_enex5;
  wire rva_out_reg_data_and_94_enex5;
  wire rva_out_reg_data_and_95_enex5;
  wire weight_port_read_out_data_and_98_enex5;
  wire rva_out_reg_data_and_96_enex5;
  wire rva_out_reg_data_and_97_enex5;
  wire rva_out_reg_data_and_98_enex5;
  wire rva_out_reg_data_and_99_enex5;
  wire rva_out_reg_data_and_100_enex5;
  wire weight_mem_write_arbxbar_xbar_for_empty_and_enex5;
  wire input_mem_banks_read_read_data_and_39_enex5;
  wire input_mem_banks_read_read_data_and_40_enex5;
  wire input_mem_banks_read_read_data_and_41_enex5;
  wire input_mem_banks_read_read_data_and_42_enex5;
  wire input_mem_banks_read_1_read_data_and_4_enex5;
  wire rva_out_reg_data_and_101_enex5;
  wire rva_out_reg_data_and_102_enex5;
  wire rva_out_reg_data_and_103_enex5;
  wire input_mem_banks_read_read_data_and_27_enex5;
  wire input_mem_banks_read_1_read_data_and_5_enex5;
  wire rva_out_reg_data_and_104_enex5;
  wire rva_out_reg_data_and_105_enex5;
  wire rva_out_reg_data_and_106_enex5;
  wire input_mem_banks_read_read_data_and_28_enex5;
  wire rva_out_reg_data_and_50_enex5;
  wire rva_out_reg_data_and_107_enex5;
  wire rva_out_reg_data_and_108_enex5;
  wire rva_out_reg_data_and_109_enex5;
  wire rva_out_reg_data_and_110_enex5;
  wire rva_out_reg_data_and_111_enex5;
  wire rva_out_reg_data_and_112_enex5;
  wire rva_out_reg_data_and_113_enex5;
  wire rva_out_reg_data_and_114_enex5;
  wire rva_out_reg_data_and_115_enex5;
  wire rva_out_reg_data_and_116_enex5;
  wire rva_out_reg_data_and_117_enex5;
  wire rva_out_reg_data_and_118_enex5;
  wire rva_out_reg_data_and_119_enex5;
  wire rva_out_reg_data_and_120_enex5;
  wire rva_out_reg_data_and_78_enex5;
  wire rva_out_reg_data_and_121_enex5;
  wire rva_out_reg_data_and_122_enex5;
  wire rva_out_reg_data_and_123_enex5;
  wire rva_out_reg_data_and_124_enex5;
  wire rva_out_reg_data_and_125_enex5;
  wire weight_port_read_out_data_and_99_enex5;
  wire weight_port_read_out_data_and_100_enex5;
  wire rva_out_reg_data_and_126_enex5;
  wire rva_out_reg_data_and_127_enex5;
  wire rva_out_reg_data_and_128_enex5;
  wire rva_out_reg_data_and_129_enex5;
  wire rva_out_reg_data_and_130_enex5;
  wire rva_out_reg_data_and_131_enex5;
  wire rva_out_reg_data_and_132_enex5;
  wire weight_port_read_out_data_and_101_enex5;
  wire weight_port_read_out_data_and_102_enex5;
  wire rva_out_reg_data_and_133_enex5;
  wire rva_out_reg_data_and_134_enex5;
  wire rva_out_reg_data_and_135_enex5;
  wire weight_port_read_out_data_and_103_enex5;
  wire weight_port_read_out_data_and_104_enex5;
  wire weight_port_read_out_data_and_105_enex5;
  wire weight_port_read_out_data_and_106_enex5;
  wire rva_out_reg_data_and_136_enex5;
  wire rva_out_reg_data_and_137_enex5;
  wire rva_out_reg_data_and_138_enex5;
  wire rva_out_reg_data_and_139_enex5;
  wire rva_out_reg_data_and_140_enex5;
  wire weight_port_read_out_data_and_107_enex5;
  wire weight_port_read_out_data_and_108_enex5;
  wire weight_port_read_out_data_and_109_enex5;
  wire weight_port_read_out_data_and_110_enex5;
  wire data_in_tmp_operator_2_for_and_tmp;
  wire pe_manager_base_input_and_tmp;
  wire rva_in_reg_data_and_tmp;
  wire and_1656_tmp;
  wire and_1694_tmp;
  wire and_1320_tmp;
  wire and_1654_tmp;
  wire and_1322_tmp;
  wire and_1776_tmp;
  wire and_1720_tmp;
  wire and_1504_tmp;
  wire and_1454_tmp;
  wire and_1304_tmp;
  wire and_1332_tmp;
  wire and_1422_tmp;
  wire and_1370_tmp;
  wire and_1542_tmp;
  wire and_1588_tmp;
  wire and_1592_tmp;
  wire and_1764_tmp;
  wire and_1576_tmp;
  wire and_1376_tmp;
  wire and_1718_tmp;
  wire and_1458_tmp;
  wire and_1444_tmp;
  wire and_1440_tmp;
  wire and_1760_tmp;
  wire and_1378_tmp;
  wire and_1470_tmp;
  wire and_1524_tmp;
  wire and_1302_tmp;
  wire and_1778_tmp;
  wire and_1774_tmp;
  wire and_1770_tmp;
  wire and_1468_tmp;
  wire and_1788_tmp;
  wire and_1312_tmp;
  wire and_1748_tmp;
  wire and_1706_tmp;
  wire and_1780_tmp;
  wire and_1740_tmp;
  wire and_1486_tmp;
  wire and_1562_tmp;
  wire and_1496_tmp;
  wire and_1350_tmp;
  wire and_1294_tmp;
  wire and_1316_tmp;
  wire and_1640_tmp;
  wire and_1632_tmp;
  wire and_1660_tmp;
  wire and_1286_tmp;
  wire and_1686_tmp;
  wire and_1384_tmp;
  wire and_1510_tmp;
  wire and_1556_tmp;
  wire and_1498_tmp;
  wire and_1550_tmp;
  wire and_1460_tmp;
  wire and_1388_tmp;
  wire and_1414_tmp;
  wire and_1726_tmp;
  wire and_1724_tmp;
  wire and_1464_tmp;
  wire and_1428_tmp;
  wire and_1548_tmp;
  wire and_1578_tmp;
  wire and_1494_tmp;
  wire and_1616_tmp;
  wire and_1382_tmp;
  wire and_1758_tmp;
  wire and_1704_tmp;
  wire and_1520_tmp;
  wire and_1306_tmp;
  wire and_1662_tmp;
  wire and_1666_tmp;
  wire and_1622_tmp;
  wire and_1512_tmp;
  wire and_1672_tmp;
  wire and_1420_tmp;
  wire and_1340_tmp;
  wire and_1360_tmp;
  wire and_1594_tmp;
  wire and_1394_tmp;
  wire and_1430_tmp;
  wire and_1326_tmp;
  wire and_1408_tmp;
  wire and_1358_tmp;
  wire and_1338_tmp;
  wire and_1580_tmp;
  wire and_1366_tmp;
  wire and_1492_tmp;
  wire and_1280_tmp;
  wire and_1356_tmp;
  wire and_1400_tmp;
  wire and_1552_tmp;
  wire and_1722_tmp;
  wire and_1608_tmp;
  wire and_1466_tmp;
  wire and_1786_tmp;
  wire and_1692_tmp;
  wire and_1372_tmp;
  wire and_1456_tmp;
  wire and_1734_tmp;
  wire and_1746_tmp;
  wire and_1664_tmp;
  wire and_1652_tmp;
  wire and_1368_tmp;
  wire and_1502_tmp;
  wire and_1300_tmp;
  wire and_1410_tmp;
  wire and_1308_tmp;
  wire and_1646_tmp;
  wire and_1484_tmp;
  wire and_1526_tmp;
  wire and_1642_tmp;
  wire and_1772_tmp;
  wire and_1446_tmp;
  wire and_1612_tmp;
  wire and_1574_tmp;
  wire and_1732_tmp;
  wire and_1742_tmp;
  wire and_1650_tmp;
  wire and_1784_tmp;
  wire and_1488_tmp;
  wire and_1480_tmp;
  wire and_1292_tmp;
  wire and_1288_tmp;
  wire and_1680_tmp;
  wire and_1750_tmp;
  wire and_1668_tmp;
  wire and_1402_tmp;
  wire and_1462_tmp;
  wire and_1314_tmp;
  wire and_1348_tmp;
  wire and_1698_tmp;
  wire and_1490_tmp;
  wire and_1418_tmp;
  wire and_1530_tmp;
  wire input_mem_banks_read_read_data_and_30_tmp;
  wire and_1284_tmp;
  wire and_1472_tmp;
  wire and_1782_tmp;
  wire and_1432_tmp;
  wire and_1392_tmp;
  wire and_1712_tmp;
  wire and_1604_tmp;
  wire and_1310_tmp;
  wire and_1362_tmp;
  wire and_1716_tmp;
  wire and_1728_tmp;
  wire and_1518_tmp;
  wire and_1404_tmp;
  wire and_1736_tmp;
  wire and_1630_tmp;
  wire and_1386_tmp;
  wire and_1426_tmp;
  wire and_1438_tmp;
  wire and_1434_tmp;
  wire and_1558_tmp;
  wire and_1584_tmp;
  wire and_1626_tmp;
  wire and_1590_tmp;
  wire and_1682_tmp;
  wire and_1754_tmp;
  wire and_1412_tmp;
  wire and_1452_tmp;
  wire and_1572_tmp;
  wire and_1618_tmp;
  wire and_1282_tmp;
  wire and_1336_tmp;
  wire and_1644_tmp;
  wire and_1610_tmp;
  wire and_1344_tmp;
  wire and_1546_tmp;
  wire and_1602_tmp;
  wire and_1596_tmp;
  wire and_1380_tmp;
  wire and_1582_tmp;
  wire and_1624_tmp;
  wire and_1636_tmp;
  wire and_1638_tmp;
  wire and_1566_tmp;
  wire and_1696_tmp;
  wire and_1374_tmp;
  wire and_1598_tmp;
  wire and_1684_tmp;
  wire and_1318_tmp;
  wire and_1364_tmp;
  wire and_1752_tmp;
  wire and_1482_tmp;
  wire and_1500_tmp;
  wire and_1536_tmp;
  wire and_1478_tmp;
  wire and_1298_tmp;
  wire and_1568_tmp;
  wire and_1756_tmp;
  wire and_1670_tmp;
  wire and_1390_tmp;
  wire and_1586_tmp;
  wire and_1560_tmp;
  wire and_1768_tmp;
  wire and_1534_tmp;
  wire and_1606_tmp;
  wire and_1628_tmp;
  wire and_1416_tmp;
  wire and_1290_tmp;
  wire and_1528_tmp;
  wire and_1532_tmp;
  wire and_1442_tmp;
  wire and_1328_tmp;
  wire and_1730_tmp;
  wire and_1554_tmp;
  wire and_1544_tmp;
  wire and_1352_tmp;
  wire and_1762_tmp;
  wire and_1620_tmp;
  wire and_1710_tmp;
  wire and_1690_tmp;
  wire and_1296_tmp;
  wire and_1342_tmp;
  wire and_1450_tmp;
  wire and_1522_tmp;
  wire and_1330_tmp;
  wire and_1658_tmp;
  wire and_1676_tmp;
  wire and_1424_tmp;
  wire and_1436_tmp;
  wire and_1506_tmp;
  wire and_1540_tmp;
  wire and_1674_tmp;
  wire and_1474_tmp;
  wire and_1614_tmp;
  wire and_1570_tmp;
  wire and_1700_tmp;
  wire and_1744_tmp;
  wire and_1508_tmp;
  wire and_1708_tmp;
  wire and_1702_tmp;
  wire and_1678_tmp;
  wire and_1564_tmp;
  wire and_1648_tmp;
  wire and_1324_tmp;
  wire and_1688_tmp;
  wire and_1476_tmp;
  wire and_1354_tmp;
  wire and_1738_tmp;
  wire and_1714_tmp;
  wire and_1766_tmp;
  wire and_1600_tmp;
  wire and_1398_tmp;
  wire and_1538_tmp;
  wire and_1634_tmp;
  wire and_1516_tmp;
  wire and_1514_tmp;
  wire and_1346_tmp;
  wire and_1334_tmp;
  wire and_1448_tmp;
  wire and_1406_tmp;
  wire and_1396_tmp;
  wire and_1278_tmp;
  wire input_mem_banks_read_read_data_and_29_tmp;
  wire rva_in_reg_rw_and_5_cse;
  wire and_990_itm;
  wire and_702_itm;
  wire mux_181_itm;
  wire mux_179_itm;
  wire mux_223_itm;
  wire mux_221_itm;
  wire PECore_PushAxiRsp_if_else_mux_14_itm;
  wire PECore_PushAxiRsp_if_else_mux_15_itm;
  wire PECore_PushAxiRsp_if_else_mux_16_itm;
  wire and_709_cse;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27;
  wire mux_101_nl;
  wire or_705_nl;
  wire mux_100_nl;
  wire nand_2_nl;
  wire mux_105_nl;
  wire or_347_nl;
  wire mux_104_nl;
  wire nand_4_nl;
  wire mux_107_nl;
  wire or_353_nl;
  wire or_351_nl;
  wire mux_109_nl;
  wire or_360_nl;
  wire or_357_nl;
  wire mux_112_nl;
  wire mux_111_nl;
  wire or_367_nl;
  wire or_365_nl;
  wire mux_118_nl;
  wire mux_117_nl;
  wire mux_116_nl;
  wire or_375_nl;
  wire mux_115_nl;
  wire or_370_nl;
  wire mux_122_nl;
  wire mux_121_nl;
  wire or_383_nl;
  wire mux_120_nl;
  wire or_381_nl;
  wire mux_128_nl;
  wire mux_127_nl;
  wire mux_126_nl;
  wire or_391_nl;
  wire mux_125_nl;
  wire or_386_nl;
  wire mux_141_nl;
  wire mux_140_nl;
  wire mux_139_nl;
  wire mux_138_nl;
  wire mux_137_nl;
  wire mux_924_nl;
  wire and_708_nl;
  wire mux_133_nl;
  wire mux_322_nl;
  wire mux_136_nl;
  wire mux_135_nl;
  wire mux_134_nl;
  wire mux_925_nl;
  wire mux_926_nl;
  wire or_218_nl;
  wire or_217_nl;
  wire or_216_nl;
  wire or_215_nl;
  wire[26:0] PECore_RunScale_if_for_3_scaled_val_mul_1_nl;
  wire or_418_nl;
  wire mux_6_nl;
  wire mux_5_nl;
  wire nor_296_nl;
  wire nor_297_nl;
  wire mux_8_nl;
  wire mux_7_nl;
  wire or_12_nl;
  wire or_11_nl;
  wire or_10_nl;
  wire mux_9_nl;
  wire mux_13_nl;
  wire mux_12_nl;
  wire mux_11_nl;
  wire mux_10_nl;
  wire or_25_nl;
  wire or_19_nl;
  wire or_17_nl;
  wire or_15_nl;
  wire or_13_nl;
  wire mux_339_nl;
  wire weight_mem_run_3_for_5_and_100_nl;
  wire mux_350_nl;
  wire mux_349_nl;
  wire weight_mem_run_3_for_5_and_81_nl;
  wire weight_mem_run_3_for_5_and_7_nl;
  wire mux_31_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_20_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_76_nl;
  wire mux_32_nl;
  wire nor_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_72_nl;
  wire mux_33_nl;
  wire nor_298_nl;
  wire or_69_nl;
  wire mux_35_nl;
  wire mux_34_nl;
  wire or_76_nl;
  wire or_74_nl;
  wire or_71_nl;
  wire mux_37_nl;
  wire mux_36_nl;
  wire nor_303_nl;
  wire or_78_nl;
  wire or_77_nl;
  wire mux_38_nl;
  wire mux_360_nl;
  wire mux_359_nl;
  wire nor_700_nl;
  wire nor_701_nl;
  wire[10:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl;
  wire[3:0] PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl;
  wire and_600_nl;
  wire[3:0] operator_4_false_acc_nl;
  wire[4:0] nl_operator_4_false_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_7_nl;
  wire mux_361_nl;
  wire nor_712_nl;
  wire nand_241_nl;
  wire mux_362_nl;
  wire nor_713_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_and_1_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_mux1h_15_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_nor_8_nl;
  wire[18:0] ProductSum_for_acc_21_nl;
  wire[19:0] nl_ProductSum_for_acc_21_nl;
  wire[18:0] ProductSum_for_acc_23_nl;
  wire[19:0] nl_ProductSum_for_acc_23_nl;
  wire PECore_UpdateFSM_switch_lp_not_19_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_129_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_101_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_115_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_122_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_94_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_108_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_130_nl;
  wire[7:0] mux1h_1_nl;
  wire and_922_nl;
  wire and_923_nl;
  wire and_924_nl;
  wire not_2217_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_123_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_109_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_131_nl;
  wire[7:0] mux_321_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_or_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_mux1h_17_nl;
  wire and_610_nl;
  wire and_612_nl;
  wire and_616_nl;
  wire and_620_nl;
  wire and_621_nl;
  wire and_613_nl;
  wire or_715_nl;
  wire nor_425_nl;
  wire mux_307_nl;
  wire mux_68_nl;
  wire mux_67_nl;
  wire mux_66_nl;
  wire mux_65_nl;
  wire mux_64_nl;
  wire mux_63_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_124_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_110_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_132_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_125_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_111_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_133_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_126_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_112_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_127_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_113_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_128_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_114_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_78_nl;
  wire mux_71_nl;
  wire or_244_nl;
  wire and_236_nl;
  wire nor_31_nl;
  wire mux_73_nl;
  wire mux_72_nl;
  wire nand_36_nl;
  wire nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_13_nl;
  wire or_248_nl;
  wire or_247_nl;
  wire or_245_nl;
  wire mux_74_nl;
  wire or_251_nl;
  wire and_238_nl;
  wire nor_32_nl;
  wire mux_75_nl;
  wire or_254_nl;
  wire and_239_nl;
  wire nor_33_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_19_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_nl;
  wire mux_76_nl;
  wire[26:0] PECore_RunScale_if_for_1_scaled_val_mul_1_nl;
  wire[26:0] PECore_RunScale_if_for_2_scaled_val_mul_1_nl;
  wire[26:0] PECore_RunScale_if_for_4_scaled_val_mul_1_nl;
  wire[26:0] PECore_RunScale_if_for_5_scaled_val_mul_1_nl;
  wire[26:0] PECore_RunScale_if_for_6_scaled_val_mul_1_nl;
  wire[26:0] PECore_RunScale_if_for_7_scaled_val_mul_1_nl;
  wire[26:0] PECore_RunScale_if_for_8_scaled_val_mul_1_nl;
  wire mux_78_nl;
  wire mux_77_nl;
  wire nor_307_nl;
  wire[18:0] ProductSum_for_acc_nl;
  wire[19:0] nl_ProductSum_for_acc_nl;
  wire[18:0] ProductSum_for_acc_36_nl;
  wire[19:0] nl_ProductSum_for_acc_36_nl;
  wire[18:0] ProductSum_for_acc_37_nl;
  wire[19:0] nl_ProductSum_for_acc_37_nl;
  wire PECore_UpdateFSM_switch_lp_not_32_nl;
  wire[18:0] ProductSum_for_acc_33_nl;
  wire[19:0] nl_ProductSum_for_acc_33_nl;
  wire[18:0] ProductSum_for_acc_34_nl;
  wire[19:0] nl_ProductSum_for_acc_34_nl;
  wire[18:0] ProductSum_for_acc_35_nl;
  wire[19:0] nl_ProductSum_for_acc_35_nl;
  wire PECore_UpdateFSM_switch_lp_not_21_nl;
  wire[18:0] ProductSum_for_acc_30_nl;
  wire[19:0] nl_ProductSum_for_acc_30_nl;
  wire[18:0] ProductSum_for_acc_31_nl;
  wire[19:0] nl_ProductSum_for_acc_31_nl;
  wire[18:0] ProductSum_for_acc_32_nl;
  wire[19:0] nl_ProductSum_for_acc_32_nl;
  wire PECore_UpdateFSM_switch_lp_not_33_nl;
  wire[18:0] ProductSum_for_acc_27_nl;
  wire[19:0] nl_ProductSum_for_acc_27_nl;
  wire[18:0] ProductSum_for_acc_28_nl;
  wire[19:0] nl_ProductSum_for_acc_28_nl;
  wire[18:0] ProductSum_for_acc_29_nl;
  wire[19:0] nl_ProductSum_for_acc_29_nl;
  wire PECore_UpdateFSM_switch_lp_not_37_nl;
  wire[18:0] ProductSum_for_acc_24_nl;
  wire[19:0] nl_ProductSum_for_acc_24_nl;
  wire[18:0] ProductSum_for_acc_25_nl;
  wire[19:0] nl_ProductSum_for_acc_25_nl;
  wire[18:0] ProductSum_for_acc_26_nl;
  wire[19:0] nl_ProductSum_for_acc_26_nl;
  wire PECore_UpdateFSM_switch_lp_not_34_nl;
  wire[18:0] ProductSum_for_acc_18_nl;
  wire[19:0] nl_ProductSum_for_acc_18_nl;
  wire[18:0] ProductSum_for_acc_19_nl;
  wire[19:0] nl_ProductSum_for_acc_19_nl;
  wire[18:0] ProductSum_for_acc_20_nl;
  wire[19:0] nl_ProductSum_for_acc_20_nl;
  wire PECore_UpdateFSM_switch_lp_not_35_nl;
  wire[18:0] ProductSum_for_acc_15_nl;
  wire[19:0] nl_ProductSum_for_acc_15_nl;
  wire[18:0] ProductSum_for_acc_16_nl;
  wire[19:0] nl_ProductSum_for_acc_16_nl;
  wire[18:0] ProductSum_for_acc_17_nl;
  wire[19:0] nl_ProductSum_for_acc_17_nl;
  wire PECore_UpdateFSM_switch_lp_not_36_nl;
  wire mux_79_nl;
  wire and_712_nl;
  wire mux_80_nl;
  wire nor_308_nl;
  wire[63:0] input_mem_banks_read_1_for_mux_4_nl;
  wire and_633_nl;
  wire nor_744_nl;
  wire nor_776_nl;
  wire nor_777_nl;
  wire or_977_nl;
  wire or_975_nl;
  wire or_1015_nl;
  wire or_1013_nl;
  wire or_1054_nl;
  wire or_1052_nl;
  wire nor_816_nl;
  wire nor_817_nl;
  wire mux_89_nl;
  wire mux_88_nl;
  wire mux_87_nl;
  wire mux_86_nl;
  wire or_317_nl;
  wire or_315_nl;
  wire or_314_nl;
  wire or_313_nl;
  wire or_312_nl;
  wire or_305_nl;
  wire weight_port_read_out_data_mux_71_nl;
  wire mux_70_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_135_nl;
  wire and_639_nl;
  wire nor_418_nl;
  wire[14:0] while_if_while_if_and_2_nl;
  wire or_492_nl;
  wire mux_90_nl;
  wire mux_92_nl;
  wire mux_91_nl;
  wire mux_93_nl;
  wire mux_95_nl;
  wire mux_94_nl;
  wire and_404_nl;
  wire or_323_nl;
  wire nor_314_nl;
  wire mux_96_nl;
  wire nor_284_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_6_nl;
  wire[63:0] input_mem_banks_bank_a_mux_1_nl;
  wire[63:0] input_mem_banks_bank_a_mux_3_nl;
  wire[63:0] input_mem_banks_bank_a_mux_5_nl;
  wire[63:0] input_mem_banks_bank_a_mux_7_nl;
  wire[63:0] input_mem_banks_bank_a_mux_9_nl;
  wire[63:0] input_mem_banks_bank_a_mux_11_nl;
  wire[63:0] input_mem_banks_bank_a_mux_13_nl;
  wire[63:0] input_mem_banks_bank_a_mux_15_nl;
  wire[63:0] input_mem_banks_bank_a_mux_17_nl;
  wire[63:0] input_mem_banks_bank_a_mux_19_nl;
  wire[63:0] input_mem_banks_bank_a_mux_21_nl;
  wire[63:0] input_mem_banks_bank_a_mux_23_nl;
  wire[63:0] input_mem_banks_bank_a_mux_25_nl;
  wire[63:0] input_mem_banks_bank_a_mux_27_nl;
  wire[63:0] input_mem_banks_bank_a_mux_29_nl;
  wire[63:0] input_mem_banks_bank_a_mux_31_nl;
  wire[63:0] input_mem_banks_bank_a_mux_33_nl;
  wire[63:0] input_mem_banks_bank_a_mux_35_nl;
  wire[63:0] input_mem_banks_bank_a_mux_37_nl;
  wire[63:0] input_mem_banks_bank_a_mux_39_nl;
  wire[63:0] input_mem_banks_bank_a_mux_41_nl;
  wire[63:0] input_mem_banks_bank_a_mux_43_nl;
  wire[63:0] input_mem_banks_bank_a_mux_45_nl;
  wire[63:0] input_mem_banks_bank_a_mux_47_nl;
  wire[63:0] input_mem_banks_bank_a_mux_49_nl;
  wire[63:0] input_mem_banks_bank_a_mux_51_nl;
  wire[63:0] input_mem_banks_bank_a_mux_53_nl;
  wire[63:0] input_mem_banks_bank_a_mux_55_nl;
  wire[63:0] input_mem_banks_bank_a_mux_57_nl;
  wire[63:0] input_mem_banks_bank_a_mux_59_nl;
  wire[63:0] input_mem_banks_bank_a_mux_61_nl;
  wire[63:0] input_mem_banks_bank_a_mux_63_nl;
  wire[63:0] input_mem_banks_bank_a_mux_65_nl;
  wire[63:0] input_mem_banks_bank_a_mux_67_nl;
  wire[63:0] input_mem_banks_bank_a_mux_69_nl;
  wire[63:0] input_mem_banks_bank_a_mux_71_nl;
  wire[63:0] input_mem_banks_bank_a_mux_73_nl;
  wire[63:0] input_mem_banks_bank_a_mux_75_nl;
  wire[63:0] input_mem_banks_bank_a_mux_77_nl;
  wire[63:0] input_mem_banks_bank_a_mux_79_nl;
  wire[63:0] input_mem_banks_bank_a_mux_81_nl;
  wire[63:0] input_mem_banks_bank_a_mux_83_nl;
  wire[63:0] input_mem_banks_bank_a_mux_85_nl;
  wire[63:0] input_mem_banks_bank_a_mux_87_nl;
  wire[63:0] input_mem_banks_bank_a_mux_89_nl;
  wire[63:0] input_mem_banks_bank_a_mux_91_nl;
  wire[63:0] input_mem_banks_bank_a_mux_93_nl;
  wire[63:0] input_mem_banks_bank_a_mux_95_nl;
  wire[63:0] input_mem_banks_bank_a_mux_97_nl;
  wire[63:0] input_mem_banks_bank_a_mux_99_nl;
  wire[63:0] input_mem_banks_bank_a_mux_101_nl;
  wire[63:0] input_mem_banks_bank_a_mux_103_nl;
  wire[63:0] input_mem_banks_bank_a_mux_105_nl;
  wire[63:0] input_mem_banks_bank_a_mux_107_nl;
  wire[63:0] input_mem_banks_bank_a_mux_109_nl;
  wire[63:0] input_mem_banks_bank_a_mux_111_nl;
  wire[63:0] input_mem_banks_bank_a_mux_113_nl;
  wire[63:0] input_mem_banks_bank_a_mux_115_nl;
  wire[63:0] input_mem_banks_bank_a_mux_117_nl;
  wire[63:0] input_mem_banks_bank_a_mux_119_nl;
  wire[63:0] input_mem_banks_bank_a_mux_121_nl;
  wire[63:0] input_mem_banks_bank_a_mux_123_nl;
  wire[63:0] input_mem_banks_bank_a_mux_125_nl;
  wire[63:0] input_mem_banks_bank_a_mux_127_nl;
  wire[63:0] input_mem_banks_bank_a_mux_129_nl;
  wire[63:0] input_mem_banks_bank_a_mux_131_nl;
  wire[63:0] input_mem_banks_bank_a_mux_133_nl;
  wire[63:0] input_mem_banks_bank_a_mux_135_nl;
  wire[63:0] input_mem_banks_bank_a_mux_137_nl;
  wire[63:0] input_mem_banks_bank_a_mux_139_nl;
  wire[63:0] input_mem_banks_bank_a_mux_141_nl;
  wire[63:0] input_mem_banks_bank_a_mux_143_nl;
  wire[63:0] input_mem_banks_bank_a_mux_145_nl;
  wire[63:0] input_mem_banks_bank_a_mux_147_nl;
  wire[63:0] input_mem_banks_bank_a_mux_149_nl;
  wire[63:0] input_mem_banks_bank_a_mux_151_nl;
  wire[63:0] input_mem_banks_bank_a_mux_153_nl;
  wire[63:0] input_mem_banks_bank_a_mux_155_nl;
  wire[63:0] input_mem_banks_bank_a_mux_157_nl;
  wire[63:0] input_mem_banks_bank_a_mux_159_nl;
  wire[63:0] input_mem_banks_bank_a_mux_161_nl;
  wire[63:0] input_mem_banks_bank_a_mux_163_nl;
  wire[63:0] input_mem_banks_bank_a_mux_165_nl;
  wire[63:0] input_mem_banks_bank_a_mux_167_nl;
  wire[63:0] input_mem_banks_bank_a_mux_169_nl;
  wire[63:0] input_mem_banks_bank_a_mux_171_nl;
  wire[63:0] input_mem_banks_bank_a_mux_173_nl;
  wire[63:0] input_mem_banks_bank_a_mux_175_nl;
  wire[63:0] input_mem_banks_bank_a_mux_177_nl;
  wire[63:0] input_mem_banks_bank_a_mux_179_nl;
  wire[63:0] input_mem_banks_bank_a_mux_181_nl;
  wire[63:0] input_mem_banks_bank_a_mux_183_nl;
  wire[63:0] input_mem_banks_bank_a_mux_185_nl;
  wire[63:0] input_mem_banks_bank_a_mux_187_nl;
  wire[63:0] input_mem_banks_bank_a_mux_189_nl;
  wire[63:0] input_mem_banks_bank_a_mux_191_nl;
  wire[63:0] input_mem_banks_bank_a_mux_193_nl;
  wire[63:0] input_mem_banks_bank_a_mux_195_nl;
  wire[63:0] input_mem_banks_bank_a_mux_197_nl;
  wire[63:0] input_mem_banks_bank_a_mux_199_nl;
  wire[63:0] input_mem_banks_bank_a_mux_201_nl;
  wire[63:0] input_mem_banks_bank_a_mux_203_nl;
  wire[63:0] input_mem_banks_bank_a_mux_205_nl;
  wire[63:0] input_mem_banks_bank_a_mux_207_nl;
  wire[63:0] input_mem_banks_bank_a_mux_209_nl;
  wire[63:0] input_mem_banks_bank_a_mux_211_nl;
  wire[63:0] input_mem_banks_bank_a_mux_213_nl;
  wire[63:0] input_mem_banks_bank_a_mux_215_nl;
  wire[63:0] input_mem_banks_bank_a_mux_217_nl;
  wire[63:0] input_mem_banks_bank_a_mux_219_nl;
  wire[63:0] input_mem_banks_bank_a_mux_221_nl;
  wire[63:0] input_mem_banks_bank_a_mux_223_nl;
  wire[63:0] input_mem_banks_bank_a_mux_225_nl;
  wire[63:0] input_mem_banks_bank_a_mux_227_nl;
  wire[63:0] input_mem_banks_bank_a_mux_229_nl;
  wire[63:0] input_mem_banks_bank_a_mux_231_nl;
  wire[63:0] input_mem_banks_bank_a_mux_233_nl;
  wire[63:0] input_mem_banks_bank_a_mux_235_nl;
  wire[63:0] input_mem_banks_bank_a_mux_237_nl;
  wire[63:0] input_mem_banks_bank_a_mux_239_nl;
  wire[63:0] input_mem_banks_bank_a_mux_241_nl;
  wire[63:0] input_mem_banks_bank_a_mux_243_nl;
  wire[63:0] input_mem_banks_bank_a_mux_245_nl;
  wire[63:0] input_mem_banks_bank_a_mux_247_nl;
  wire[63:0] input_mem_banks_bank_a_mux_249_nl;
  wire[63:0] input_mem_banks_bank_a_mux_251_nl;
  wire[63:0] input_mem_banks_bank_a_mux_253_nl;
  wire[63:0] input_mem_banks_bank_a_mux_255_nl;
  wire[63:0] input_mem_banks_bank_a_mux_257_nl;
  wire[63:0] input_mem_banks_bank_a_mux_259_nl;
  wire[63:0] input_mem_banks_bank_a_mux_261_nl;
  wire[63:0] input_mem_banks_bank_a_mux_263_nl;
  wire[63:0] input_mem_banks_bank_a_mux_265_nl;
  wire[63:0] input_mem_banks_bank_a_mux_267_nl;
  wire[63:0] input_mem_banks_bank_a_mux_269_nl;
  wire[63:0] input_mem_banks_bank_a_mux_271_nl;
  wire[63:0] input_mem_banks_bank_a_mux_273_nl;
  wire[63:0] input_mem_banks_bank_a_mux_275_nl;
  wire[63:0] input_mem_banks_bank_a_mux_277_nl;
  wire[63:0] input_mem_banks_bank_a_mux_279_nl;
  wire[63:0] input_mem_banks_bank_a_mux_281_nl;
  wire[63:0] input_mem_banks_bank_a_mux_283_nl;
  wire[63:0] input_mem_banks_bank_a_mux_285_nl;
  wire[63:0] input_mem_banks_bank_a_mux_287_nl;
  wire[63:0] input_mem_banks_bank_a_mux_289_nl;
  wire[63:0] input_mem_banks_bank_a_mux_291_nl;
  wire[63:0] input_mem_banks_bank_a_mux_293_nl;
  wire[63:0] input_mem_banks_bank_a_mux_295_nl;
  wire[63:0] input_mem_banks_bank_a_mux_297_nl;
  wire[63:0] input_mem_banks_bank_a_mux_299_nl;
  wire[63:0] input_mem_banks_bank_a_mux_301_nl;
  wire[63:0] input_mem_banks_bank_a_mux_303_nl;
  wire[63:0] input_mem_banks_bank_a_mux_305_nl;
  wire[63:0] input_mem_banks_bank_a_mux_307_nl;
  wire[63:0] input_mem_banks_bank_a_mux_309_nl;
  wire[63:0] input_mem_banks_bank_a_mux_311_nl;
  wire[63:0] input_mem_banks_bank_a_mux_313_nl;
  wire[63:0] input_mem_banks_bank_a_mux_315_nl;
  wire[63:0] input_mem_banks_bank_a_mux_317_nl;
  wire[63:0] input_mem_banks_bank_a_mux_319_nl;
  wire[63:0] input_mem_banks_bank_a_mux_321_nl;
  wire[63:0] input_mem_banks_bank_a_mux_323_nl;
  wire[63:0] input_mem_banks_bank_a_mux_325_nl;
  wire[63:0] input_mem_banks_bank_a_mux_327_nl;
  wire[63:0] input_mem_banks_bank_a_mux_329_nl;
  wire[63:0] input_mem_banks_bank_a_mux_331_nl;
  wire[63:0] input_mem_banks_bank_a_mux_333_nl;
  wire[63:0] input_mem_banks_bank_a_mux_335_nl;
  wire[63:0] input_mem_banks_bank_a_mux_337_nl;
  wire[63:0] input_mem_banks_bank_a_mux_339_nl;
  wire[63:0] input_mem_banks_bank_a_mux_341_nl;
  wire[63:0] input_mem_banks_bank_a_mux_343_nl;
  wire[63:0] input_mem_banks_bank_a_mux_345_nl;
  wire[63:0] input_mem_banks_bank_a_mux_347_nl;
  wire[63:0] input_mem_banks_bank_a_mux_349_nl;
  wire[63:0] input_mem_banks_bank_a_mux_351_nl;
  wire[63:0] input_mem_banks_bank_a_mux_353_nl;
  wire[63:0] input_mem_banks_bank_a_mux_355_nl;
  wire[63:0] input_mem_banks_bank_a_mux_357_nl;
  wire[63:0] input_mem_banks_bank_a_mux_359_nl;
  wire[63:0] input_mem_banks_bank_a_mux_361_nl;
  wire[63:0] input_mem_banks_bank_a_mux_363_nl;
  wire[63:0] input_mem_banks_bank_a_mux_365_nl;
  wire[63:0] input_mem_banks_bank_a_mux_367_nl;
  wire[63:0] input_mem_banks_bank_a_mux_369_nl;
  wire[63:0] input_mem_banks_bank_a_mux_371_nl;
  wire[63:0] input_mem_banks_bank_a_mux_373_nl;
  wire[63:0] input_mem_banks_bank_a_mux_375_nl;
  wire[63:0] input_mem_banks_bank_a_mux_377_nl;
  wire[63:0] input_mem_banks_bank_a_mux_379_nl;
  wire[63:0] input_mem_banks_bank_a_mux_381_nl;
  wire[63:0] input_mem_banks_bank_a_mux_383_nl;
  wire[63:0] input_mem_banks_bank_a_mux_385_nl;
  wire[63:0] input_mem_banks_bank_a_mux_387_nl;
  wire[63:0] input_mem_banks_bank_a_mux_389_nl;
  wire[63:0] input_mem_banks_bank_a_mux_391_nl;
  wire[63:0] input_mem_banks_bank_a_mux_393_nl;
  wire[63:0] input_mem_banks_bank_a_mux_395_nl;
  wire[63:0] input_mem_banks_bank_a_mux_397_nl;
  wire[63:0] input_mem_banks_bank_a_mux_399_nl;
  wire[63:0] input_mem_banks_bank_a_mux_401_nl;
  wire[63:0] input_mem_banks_bank_a_mux_403_nl;
  wire[63:0] input_mem_banks_bank_a_mux_405_nl;
  wire[63:0] input_mem_banks_bank_a_mux_407_nl;
  wire[63:0] input_mem_banks_bank_a_mux_409_nl;
  wire[63:0] input_mem_banks_bank_a_mux_411_nl;
  wire[63:0] input_mem_banks_bank_a_mux_413_nl;
  wire[63:0] input_mem_banks_bank_a_mux_415_nl;
  wire[63:0] input_mem_banks_bank_a_mux_417_nl;
  wire[63:0] input_mem_banks_bank_a_mux_419_nl;
  wire[63:0] input_mem_banks_bank_a_mux_421_nl;
  wire[63:0] input_mem_banks_bank_a_mux_423_nl;
  wire[63:0] input_mem_banks_bank_a_mux_425_nl;
  wire[63:0] input_mem_banks_bank_a_mux_427_nl;
  wire[63:0] input_mem_banks_bank_a_mux_429_nl;
  wire[63:0] input_mem_banks_bank_a_mux_431_nl;
  wire[63:0] input_mem_banks_bank_a_mux_433_nl;
  wire[63:0] input_mem_banks_bank_a_mux_435_nl;
  wire[63:0] input_mem_banks_bank_a_mux_437_nl;
  wire[63:0] input_mem_banks_bank_a_mux_439_nl;
  wire[63:0] input_mem_banks_bank_a_mux_441_nl;
  wire[63:0] input_mem_banks_bank_a_mux_443_nl;
  wire[63:0] input_mem_banks_bank_a_mux_445_nl;
  wire[63:0] input_mem_banks_bank_a_mux_447_nl;
  wire[63:0] input_mem_banks_bank_a_mux_449_nl;
  wire[63:0] input_mem_banks_bank_a_mux_451_nl;
  wire[63:0] input_mem_banks_bank_a_mux_453_nl;
  wire[63:0] input_mem_banks_bank_a_mux_455_nl;
  wire[63:0] input_mem_banks_bank_a_mux_457_nl;
  wire[63:0] input_mem_banks_bank_a_mux_459_nl;
  wire[63:0] input_mem_banks_bank_a_mux_461_nl;
  wire[63:0] input_mem_banks_bank_a_mux_463_nl;
  wire[63:0] input_mem_banks_bank_a_mux_465_nl;
  wire[63:0] input_mem_banks_bank_a_mux_467_nl;
  wire[63:0] input_mem_banks_bank_a_mux_469_nl;
  wire[63:0] input_mem_banks_bank_a_mux_471_nl;
  wire[63:0] input_mem_banks_bank_a_mux_473_nl;
  wire[63:0] input_mem_banks_bank_a_mux_475_nl;
  wire[63:0] input_mem_banks_bank_a_mux_477_nl;
  wire[63:0] input_mem_banks_bank_a_mux_479_nl;
  wire[63:0] input_mem_banks_bank_a_mux_481_nl;
  wire[63:0] input_mem_banks_bank_a_mux_483_nl;
  wire[63:0] input_mem_banks_bank_a_mux_485_nl;
  wire[63:0] input_mem_banks_bank_a_mux_487_nl;
  wire[63:0] input_mem_banks_bank_a_mux_489_nl;
  wire[63:0] input_mem_banks_bank_a_mux_491_nl;
  wire[63:0] input_mem_banks_bank_a_mux_493_nl;
  wire[63:0] input_mem_banks_bank_a_mux_495_nl;
  wire[63:0] input_mem_banks_bank_a_mux_497_nl;
  wire[63:0] input_mem_banks_bank_a_mux_499_nl;
  wire[63:0] input_mem_banks_bank_a_mux_501_nl;
  wire[63:0] input_mem_banks_bank_a_mux_503_nl;
  wire[63:0] input_mem_banks_bank_a_mux_505_nl;
  wire[63:0] input_mem_banks_bank_a_mux_507_nl;
  wire[63:0] input_mem_banks_bank_a_mux_509_nl;
  wire[63:0] input_mem_banks_bank_a_mux_511_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_74_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_76_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_77_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_79_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_92_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_95_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl;
  wire[14:0] PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_nl;
  wire[14:0] nl_operator_15_false_acc_nl;
  wire[14:0] PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[12:0] operator_15_false_acc_1_nl;
  wire[13:0] nl_operator_15_false_acc_1_nl;
  wire[14:0] PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_2_nl;
  wire[14:0] nl_operator_15_false_acc_2_nl;
  wire[14:0] PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl;
  wire and_628_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl;
  wire[7:0] pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl;
  wire[7:0] operator_8_false_acc_nl;
  wire[8:0] nl_operator_8_false_acc_nl;
  wire pe_config_UpdateInputCounter_not_nl;
  wire pe_config_input_counter_nand_nl;
  wire while_and_4_nl;
  wire[7:0] pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl;
  wire[7:0] operator_8_false_1_acc_nl;
  wire[8:0] nl_operator_8_false_1_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_9_nl;
  wire pe_config_output_counter_nand_nl;
  wire while_and_63_nl;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl;
  wire while_if_or_nl;
  wire while_if_and_4_nl;
  wire[15:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_nl;
  wire PECore_UpdateFSM_switch_lp_not_16_nl;
  wire or_452_nl;
  wire[15:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_nl;
  wire PECore_UpdateFSM_switch_lp_not_26_nl;
  wire[15:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_nl;
  wire PECore_UpdateFSM_switch_lp_not_27_nl;
  wire[15:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_nl;
  wire PECore_UpdateFSM_switch_lp_not_28_nl;
  wire[15:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_11_nl;
  wire PECore_UpdateFSM_switch_lp_not_29_nl;
  wire[15:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_10_nl;
  wire PECore_UpdateFSM_switch_lp_not_30_nl;
  wire[15:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_9_nl;
  wire PECore_UpdateFSM_switch_lp_not_31_nl;
  wire[15:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl;
  wire PECore_UpdateFSM_switch_lp_not_25_nl;
  wire while_or_2_nl;
  wire while_and_100_nl;
  wire while_and_101_nl;
  wire while_or_3_nl;
  wire while_and_104_nl;
  wire while_and_105_nl;
  wire while_or_4_nl;
  wire while_and_108_nl;
  wire while_and_109_nl;
  wire while_or_5_nl;
  wire while_and_112_nl;
  wire while_and_113_nl;
  wire while_or_6_nl;
  wire while_and_116_nl;
  wire while_and_117_nl;
  wire while_or_7_nl;
  wire while_and_120_nl;
  wire while_and_121_nl;
  wire while_or_8_nl;
  wire while_and_124_nl;
  wire while_and_125_nl;
  wire while_or_9_nl;
  wire while_and_128_nl;
  wire while_and_129_nl;
  wire while_or_10_nl;
  wire while_and_132_nl;
  wire while_and_133_nl;
  wire while_or_11_nl;
  wire while_and_136_nl;
  wire while_and_137_nl;
  wire while_or_12_nl;
  wire while_and_140_nl;
  wire while_and_141_nl;
  wire while_or_13_nl;
  wire while_and_144_nl;
  wire while_and_145_nl;
  wire while_or_14_nl;
  wire while_and_148_nl;
  wire while_and_149_nl;
  wire while_or_15_nl;
  wire while_and_152_nl;
  wire while_and_153_nl;
  wire while_or_16_nl;
  wire while_and_156_nl;
  wire while_and_157_nl;
  wire while_or_17_nl;
  wire while_and_160_nl;
  wire while_and_161_nl;
  wire while_or_18_nl;
  wire while_and_164_nl;
  wire while_and_165_nl;
  wire while_or_19_nl;
  wire while_and_168_nl;
  wire while_and_169_nl;
  wire while_or_20_nl;
  wire while_and_172_nl;
  wire while_and_173_nl;
  wire while_or_21_nl;
  wire while_and_176_nl;
  wire while_and_177_nl;
  wire while_or_22_nl;
  wire while_and_180_nl;
  wire while_and_181_nl;
  wire while_or_23_nl;
  wire while_and_184_nl;
  wire while_and_185_nl;
  wire while_or_24_nl;
  wire while_and_188_nl;
  wire while_and_189_nl;
  wire while_or_25_nl;
  wire while_and_192_nl;
  wire while_and_193_nl;
  wire while_or_26_nl;
  wire while_and_196_nl;
  wire while_and_197_nl;
  wire while_or_27_nl;
  wire while_and_200_nl;
  wire while_and_201_nl;
  wire while_or_28_nl;
  wire while_and_204_nl;
  wire while_and_205_nl;
  wire while_or_29_nl;
  wire while_and_208_nl;
  wire while_and_209_nl;
  wire while_or_30_nl;
  wire while_and_212_nl;
  wire while_and_213_nl;
  wire while_or_31_nl;
  wire while_and_216_nl;
  wire while_and_217_nl;
  wire while_or_32_nl;
  wire while_and_220_nl;
  wire while_and_221_nl;
  wire while_or_33_nl;
  wire while_and_224_nl;
  wire while_and_225_nl;
  wire while_or_34_nl;
  wire while_and_228_nl;
  wire while_and_229_nl;
  wire while_or_35_nl;
  wire while_and_232_nl;
  wire while_and_233_nl;
  wire while_or_36_nl;
  wire while_and_236_nl;
  wire while_and_237_nl;
  wire while_or_37_nl;
  wire while_and_240_nl;
  wire while_and_241_nl;
  wire while_or_38_nl;
  wire while_and_244_nl;
  wire while_and_245_nl;
  wire while_or_39_nl;
  wire while_and_248_nl;
  wire while_and_249_nl;
  wire while_or_40_nl;
  wire while_and_252_nl;
  wire while_and_253_nl;
  wire while_or_41_nl;
  wire while_and_256_nl;
  wire while_and_257_nl;
  wire while_or_42_nl;
  wire while_and_260_nl;
  wire while_and_261_nl;
  wire while_or_43_nl;
  wire while_and_264_nl;
  wire while_and_265_nl;
  wire while_or_44_nl;
  wire while_and_268_nl;
  wire while_and_269_nl;
  wire while_or_45_nl;
  wire while_and_272_nl;
  wire while_and_273_nl;
  wire while_or_46_nl;
  wire while_and_276_nl;
  wire while_and_277_nl;
  wire while_or_47_nl;
  wire while_and_280_nl;
  wire while_and_281_nl;
  wire while_or_48_nl;
  wire while_and_284_nl;
  wire while_and_285_nl;
  wire while_or_49_nl;
  wire while_and_288_nl;
  wire while_and_289_nl;
  wire while_or_50_nl;
  wire while_and_292_nl;
  wire while_and_293_nl;
  wire while_or_51_nl;
  wire while_and_296_nl;
  wire while_and_297_nl;
  wire while_or_52_nl;
  wire while_and_300_nl;
  wire while_and_301_nl;
  wire while_or_53_nl;
  wire while_and_304_nl;
  wire while_and_305_nl;
  wire while_or_54_nl;
  wire while_and_308_nl;
  wire while_and_309_nl;
  wire while_or_55_nl;
  wire while_and_312_nl;
  wire while_and_313_nl;
  wire while_or_56_nl;
  wire while_and_316_nl;
  wire while_and_317_nl;
  wire while_or_57_nl;
  wire while_and_320_nl;
  wire while_and_321_nl;
  wire while_or_58_nl;
  wire while_and_324_nl;
  wire while_and_325_nl;
  wire while_or_59_nl;
  wire while_and_328_nl;
  wire while_and_329_nl;
  wire while_or_60_nl;
  wire while_and_332_nl;
  wire while_and_333_nl;
  wire while_or_61_nl;
  wire while_and_336_nl;
  wire while_and_337_nl;
  wire while_or_62_nl;
  wire while_and_340_nl;
  wire while_and_341_nl;
  wire while_or_63_nl;
  wire while_and_344_nl;
  wire while_and_345_nl;
  wire while_or_64_nl;
  wire while_and_348_nl;
  wire while_and_349_nl;
  wire while_or_65_nl;
  wire while_and_352_nl;
  wire while_and_353_nl;
  wire while_or_66_nl;
  wire while_and_356_nl;
  wire while_and_357_nl;
  wire while_or_67_nl;
  wire while_and_360_nl;
  wire while_and_361_nl;
  wire while_or_68_nl;
  wire while_and_364_nl;
  wire while_and_365_nl;
  wire while_or_69_nl;
  wire while_and_368_nl;
  wire while_and_369_nl;
  wire while_or_70_nl;
  wire while_and_372_nl;
  wire while_and_373_nl;
  wire while_or_71_nl;
  wire while_and_376_nl;
  wire while_and_377_nl;
  wire while_or_72_nl;
  wire while_and_380_nl;
  wire while_and_381_nl;
  wire while_or_73_nl;
  wire while_and_384_nl;
  wire while_and_385_nl;
  wire while_or_74_nl;
  wire while_and_388_nl;
  wire while_and_389_nl;
  wire while_or_75_nl;
  wire while_and_392_nl;
  wire while_and_393_nl;
  wire while_or_76_nl;
  wire while_and_396_nl;
  wire while_and_397_nl;
  wire while_or_77_nl;
  wire while_and_400_nl;
  wire while_and_401_nl;
  wire while_or_78_nl;
  wire while_and_404_nl;
  wire while_and_405_nl;
  wire while_or_79_nl;
  wire while_and_408_nl;
  wire while_and_409_nl;
  wire while_or_80_nl;
  wire while_and_412_nl;
  wire while_and_413_nl;
  wire while_or_81_nl;
  wire while_and_416_nl;
  wire while_and_417_nl;
  wire while_or_82_nl;
  wire while_and_420_nl;
  wire while_and_421_nl;
  wire while_or_83_nl;
  wire while_and_424_nl;
  wire while_and_425_nl;
  wire while_or_84_nl;
  wire while_and_428_nl;
  wire while_and_429_nl;
  wire while_or_85_nl;
  wire while_and_432_nl;
  wire while_and_433_nl;
  wire while_or_86_nl;
  wire while_and_436_nl;
  wire while_and_437_nl;
  wire while_or_87_nl;
  wire while_and_440_nl;
  wire while_and_441_nl;
  wire while_or_88_nl;
  wire while_and_444_nl;
  wire while_and_445_nl;
  wire while_or_89_nl;
  wire while_and_448_nl;
  wire while_and_449_nl;
  wire while_or_90_nl;
  wire while_and_452_nl;
  wire while_and_453_nl;
  wire while_or_91_nl;
  wire while_and_456_nl;
  wire while_and_457_nl;
  wire while_or_92_nl;
  wire while_and_460_nl;
  wire while_and_461_nl;
  wire while_or_93_nl;
  wire while_and_464_nl;
  wire while_and_465_nl;
  wire while_or_94_nl;
  wire while_and_468_nl;
  wire while_and_469_nl;
  wire while_or_95_nl;
  wire while_and_472_nl;
  wire while_and_473_nl;
  wire while_or_96_nl;
  wire while_and_476_nl;
  wire while_and_477_nl;
  wire while_or_97_nl;
  wire while_and_480_nl;
  wire while_and_481_nl;
  wire while_or_98_nl;
  wire while_and_484_nl;
  wire while_and_485_nl;
  wire while_or_99_nl;
  wire while_and_488_nl;
  wire while_and_489_nl;
  wire while_or_100_nl;
  wire while_and_492_nl;
  wire while_and_493_nl;
  wire while_or_101_nl;
  wire while_and_496_nl;
  wire while_and_497_nl;
  wire while_or_102_nl;
  wire while_and_500_nl;
  wire while_and_501_nl;
  wire while_or_103_nl;
  wire while_and_504_nl;
  wire while_and_505_nl;
  wire while_or_104_nl;
  wire while_and_508_nl;
  wire while_and_509_nl;
  wire while_or_105_nl;
  wire while_and_512_nl;
  wire while_and_513_nl;
  wire while_or_106_nl;
  wire while_and_516_nl;
  wire while_and_517_nl;
  wire while_or_107_nl;
  wire while_and_520_nl;
  wire while_and_521_nl;
  wire while_or_108_nl;
  wire while_and_524_nl;
  wire while_and_525_nl;
  wire while_or_109_nl;
  wire while_and_528_nl;
  wire while_and_529_nl;
  wire while_or_110_nl;
  wire while_and_532_nl;
  wire while_and_533_nl;
  wire while_or_111_nl;
  wire while_and_536_nl;
  wire while_and_537_nl;
  wire while_or_112_nl;
  wire while_and_540_nl;
  wire while_and_541_nl;
  wire while_or_113_nl;
  wire while_and_544_nl;
  wire while_and_545_nl;
  wire while_or_114_nl;
  wire while_and_548_nl;
  wire while_and_549_nl;
  wire while_or_115_nl;
  wire while_and_552_nl;
  wire while_and_553_nl;
  wire while_or_116_nl;
  wire while_and_556_nl;
  wire while_and_557_nl;
  wire while_or_117_nl;
  wire while_and_560_nl;
  wire while_and_561_nl;
  wire while_or_118_nl;
  wire while_and_564_nl;
  wire while_and_565_nl;
  wire while_or_119_nl;
  wire while_and_568_nl;
  wire while_and_569_nl;
  wire while_or_120_nl;
  wire while_and_572_nl;
  wire while_and_573_nl;
  wire while_or_121_nl;
  wire while_and_576_nl;
  wire while_and_577_nl;
  wire while_or_122_nl;
  wire while_and_580_nl;
  wire while_and_581_nl;
  wire while_or_123_nl;
  wire while_and_584_nl;
  wire while_and_585_nl;
  wire while_or_124_nl;
  wire while_and_588_nl;
  wire while_and_589_nl;
  wire while_or_125_nl;
  wire while_and_592_nl;
  wire while_and_593_nl;
  wire while_or_126_nl;
  wire while_and_596_nl;
  wire while_and_597_nl;
  wire while_or_127_nl;
  wire while_and_600_nl;
  wire while_and_601_nl;
  wire while_or_128_nl;
  wire while_and_604_nl;
  wire while_and_605_nl;
  wire while_or_129_nl;
  wire while_and_608_nl;
  wire while_and_609_nl;
  wire while_or_130_nl;
  wire while_and_612_nl;
  wire while_and_613_nl;
  wire while_or_131_nl;
  wire while_and_616_nl;
  wire while_and_617_nl;
  wire while_or_132_nl;
  wire while_and_620_nl;
  wire while_and_621_nl;
  wire while_or_133_nl;
  wire while_and_624_nl;
  wire while_and_625_nl;
  wire while_or_134_nl;
  wire while_and_628_nl;
  wire while_and_629_nl;
  wire while_or_135_nl;
  wire while_and_632_nl;
  wire while_and_633_nl;
  wire while_or_136_nl;
  wire while_and_636_nl;
  wire while_and_637_nl;
  wire while_or_137_nl;
  wire while_and_640_nl;
  wire while_and_641_nl;
  wire while_or_138_nl;
  wire while_and_644_nl;
  wire while_and_645_nl;
  wire while_or_139_nl;
  wire while_and_648_nl;
  wire while_and_649_nl;
  wire while_or_140_nl;
  wire while_and_652_nl;
  wire while_and_653_nl;
  wire while_or_141_nl;
  wire while_and_656_nl;
  wire while_and_657_nl;
  wire while_or_142_nl;
  wire while_and_660_nl;
  wire while_and_661_nl;
  wire while_or_143_nl;
  wire while_and_664_nl;
  wire while_and_665_nl;
  wire while_or_144_nl;
  wire while_and_668_nl;
  wire while_and_669_nl;
  wire while_or_145_nl;
  wire while_and_672_nl;
  wire while_and_673_nl;
  wire while_or_146_nl;
  wire while_and_676_nl;
  wire while_and_677_nl;
  wire while_or_147_nl;
  wire while_and_680_nl;
  wire while_and_681_nl;
  wire while_or_148_nl;
  wire while_and_684_nl;
  wire while_and_685_nl;
  wire while_or_149_nl;
  wire while_and_688_nl;
  wire while_and_689_nl;
  wire while_or_150_nl;
  wire while_and_692_nl;
  wire while_and_693_nl;
  wire while_or_151_nl;
  wire while_and_696_nl;
  wire while_and_697_nl;
  wire while_or_152_nl;
  wire while_and_700_nl;
  wire while_and_701_nl;
  wire while_or_153_nl;
  wire while_and_704_nl;
  wire while_and_705_nl;
  wire while_or_154_nl;
  wire while_and_708_nl;
  wire while_and_709_nl;
  wire while_or_155_nl;
  wire while_and_712_nl;
  wire while_and_713_nl;
  wire while_or_156_nl;
  wire while_and_716_nl;
  wire while_and_717_nl;
  wire while_or_157_nl;
  wire while_and_720_nl;
  wire while_and_721_nl;
  wire while_or_158_nl;
  wire while_and_724_nl;
  wire while_and_725_nl;
  wire while_or_159_nl;
  wire while_and_728_nl;
  wire while_and_729_nl;
  wire while_or_160_nl;
  wire while_and_732_nl;
  wire while_and_733_nl;
  wire while_or_161_nl;
  wire while_and_736_nl;
  wire while_and_737_nl;
  wire while_or_162_nl;
  wire while_and_740_nl;
  wire while_and_741_nl;
  wire while_or_163_nl;
  wire while_and_744_nl;
  wire while_and_745_nl;
  wire while_or_164_nl;
  wire while_and_748_nl;
  wire while_and_749_nl;
  wire while_or_165_nl;
  wire while_and_752_nl;
  wire while_and_753_nl;
  wire while_or_166_nl;
  wire while_and_756_nl;
  wire while_and_757_nl;
  wire while_or_167_nl;
  wire while_and_760_nl;
  wire while_and_761_nl;
  wire while_or_168_nl;
  wire while_and_764_nl;
  wire while_and_765_nl;
  wire while_or_169_nl;
  wire while_and_768_nl;
  wire while_and_769_nl;
  wire while_or_170_nl;
  wire while_and_772_nl;
  wire while_and_773_nl;
  wire while_or_171_nl;
  wire while_and_776_nl;
  wire while_and_777_nl;
  wire while_or_172_nl;
  wire while_and_780_nl;
  wire while_and_781_nl;
  wire while_or_173_nl;
  wire while_and_784_nl;
  wire while_and_785_nl;
  wire while_or_174_nl;
  wire while_and_788_nl;
  wire while_and_789_nl;
  wire while_or_175_nl;
  wire while_and_792_nl;
  wire while_and_793_nl;
  wire while_or_176_nl;
  wire while_and_796_nl;
  wire while_and_797_nl;
  wire while_or_177_nl;
  wire while_and_800_nl;
  wire while_and_801_nl;
  wire while_or_178_nl;
  wire while_and_804_nl;
  wire while_and_805_nl;
  wire while_or_179_nl;
  wire while_and_808_nl;
  wire while_and_809_nl;
  wire while_or_180_nl;
  wire while_and_812_nl;
  wire while_and_813_nl;
  wire while_or_181_nl;
  wire while_and_816_nl;
  wire while_and_817_nl;
  wire while_or_182_nl;
  wire while_and_820_nl;
  wire while_and_821_nl;
  wire while_or_183_nl;
  wire while_and_824_nl;
  wire while_and_825_nl;
  wire while_or_184_nl;
  wire while_and_828_nl;
  wire while_and_829_nl;
  wire while_or_185_nl;
  wire while_and_832_nl;
  wire while_and_833_nl;
  wire while_or_186_nl;
  wire while_and_836_nl;
  wire while_and_837_nl;
  wire while_or_187_nl;
  wire while_and_840_nl;
  wire while_and_841_nl;
  wire while_or_188_nl;
  wire while_and_844_nl;
  wire while_and_845_nl;
  wire while_or_189_nl;
  wire while_and_848_nl;
  wire while_and_849_nl;
  wire while_or_190_nl;
  wire while_and_852_nl;
  wire while_and_853_nl;
  wire while_or_191_nl;
  wire while_and_856_nl;
  wire while_and_857_nl;
  wire while_or_192_nl;
  wire while_and_860_nl;
  wire while_and_861_nl;
  wire while_or_193_nl;
  wire while_and_864_nl;
  wire while_and_865_nl;
  wire while_or_194_nl;
  wire while_and_868_nl;
  wire while_and_869_nl;
  wire while_or_195_nl;
  wire while_and_872_nl;
  wire while_and_873_nl;
  wire while_or_196_nl;
  wire while_and_876_nl;
  wire while_and_877_nl;
  wire while_or_197_nl;
  wire while_and_880_nl;
  wire while_and_881_nl;
  wire while_or_198_nl;
  wire while_and_884_nl;
  wire while_and_885_nl;
  wire while_or_199_nl;
  wire while_and_888_nl;
  wire while_and_889_nl;
  wire while_or_200_nl;
  wire while_and_892_nl;
  wire while_and_893_nl;
  wire while_or_201_nl;
  wire while_and_896_nl;
  wire while_and_897_nl;
  wire while_or_202_nl;
  wire while_and_900_nl;
  wire while_and_901_nl;
  wire while_or_203_nl;
  wire while_and_904_nl;
  wire while_and_905_nl;
  wire while_or_204_nl;
  wire while_and_908_nl;
  wire while_and_909_nl;
  wire while_or_205_nl;
  wire while_and_912_nl;
  wire while_and_913_nl;
  wire while_or_206_nl;
  wire while_and_916_nl;
  wire while_and_917_nl;
  wire while_or_207_nl;
  wire while_and_920_nl;
  wire while_and_921_nl;
  wire while_or_208_nl;
  wire while_and_924_nl;
  wire while_and_925_nl;
  wire while_or_209_nl;
  wire while_and_928_nl;
  wire while_and_929_nl;
  wire while_or_210_nl;
  wire while_and_932_nl;
  wire while_and_933_nl;
  wire while_or_211_nl;
  wire while_and_936_nl;
  wire while_and_937_nl;
  wire while_or_212_nl;
  wire while_and_940_nl;
  wire while_and_941_nl;
  wire while_or_213_nl;
  wire while_and_944_nl;
  wire while_and_945_nl;
  wire while_or_214_nl;
  wire while_and_948_nl;
  wire while_and_949_nl;
  wire while_or_215_nl;
  wire while_and_952_nl;
  wire while_and_953_nl;
  wire while_or_216_nl;
  wire while_and_956_nl;
  wire while_and_957_nl;
  wire while_or_217_nl;
  wire while_and_960_nl;
  wire while_and_961_nl;
  wire while_or_218_nl;
  wire while_and_964_nl;
  wire while_and_965_nl;
  wire while_or_219_nl;
  wire while_and_968_nl;
  wire while_and_969_nl;
  wire while_or_220_nl;
  wire while_and_972_nl;
  wire while_and_973_nl;
  wire while_or_221_nl;
  wire while_and_976_nl;
  wire while_and_977_nl;
  wire while_or_222_nl;
  wire while_and_980_nl;
  wire while_and_981_nl;
  wire while_or_223_nl;
  wire while_and_984_nl;
  wire while_and_985_nl;
  wire while_or_224_nl;
  wire while_and_988_nl;
  wire while_and_989_nl;
  wire while_or_225_nl;
  wire while_and_992_nl;
  wire while_and_993_nl;
  wire while_or_226_nl;
  wire while_and_996_nl;
  wire while_and_997_nl;
  wire while_or_227_nl;
  wire while_and_1000_nl;
  wire while_and_1001_nl;
  wire while_or_228_nl;
  wire while_and_1004_nl;
  wire while_and_1005_nl;
  wire while_or_229_nl;
  wire while_and_1008_nl;
  wire while_and_1009_nl;
  wire while_or_230_nl;
  wire while_and_1012_nl;
  wire while_and_1013_nl;
  wire while_or_231_nl;
  wire while_and_1016_nl;
  wire while_and_1017_nl;
  wire while_or_232_nl;
  wire while_and_1020_nl;
  wire while_and_1021_nl;
  wire while_or_233_nl;
  wire while_and_1024_nl;
  wire while_and_1025_nl;
  wire while_or_234_nl;
  wire while_and_1028_nl;
  wire while_and_1029_nl;
  wire while_or_235_nl;
  wire while_and_1032_nl;
  wire while_and_1033_nl;
  wire while_or_236_nl;
  wire while_and_1036_nl;
  wire while_and_1037_nl;
  wire while_or_237_nl;
  wire while_and_1040_nl;
  wire while_and_1041_nl;
  wire while_or_238_nl;
  wire while_and_1044_nl;
  wire while_and_1045_nl;
  wire while_or_239_nl;
  wire while_and_1048_nl;
  wire while_and_1049_nl;
  wire while_or_240_nl;
  wire while_and_1052_nl;
  wire while_and_1053_nl;
  wire while_or_241_nl;
  wire while_and_1056_nl;
  wire while_and_1057_nl;
  wire while_or_242_nl;
  wire while_and_1060_nl;
  wire while_and_1061_nl;
  wire while_or_243_nl;
  wire while_and_1064_nl;
  wire while_and_1065_nl;
  wire while_or_244_nl;
  wire while_and_1068_nl;
  wire while_and_1069_nl;
  wire while_or_245_nl;
  wire while_and_1072_nl;
  wire while_and_1073_nl;
  wire while_or_246_nl;
  wire while_and_1076_nl;
  wire while_and_1077_nl;
  wire while_or_247_nl;
  wire while_and_1080_nl;
  wire while_and_1081_nl;
  wire while_or_248_nl;
  wire while_and_1084_nl;
  wire while_and_1085_nl;
  wire while_or_249_nl;
  wire while_and_1088_nl;
  wire while_and_1089_nl;
  wire while_or_250_nl;
  wire while_and_1092_nl;
  wire while_and_1093_nl;
  wire while_or_251_nl;
  wire while_and_1096_nl;
  wire while_and_1097_nl;
  wire while_or_252_nl;
  wire while_and_1100_nl;
  wire while_and_1101_nl;
  wire while_or_253_nl;
  wire while_and_1104_nl;
  wire while_and_1105_nl;
  wire while_or_254_nl;
  wire while_and_1108_nl;
  wire while_and_1109_nl;
  wire while_or_255_nl;
  wire while_and_1112_nl;
  wire while_and_1113_nl;
  wire while_or_256_nl;
  wire while_and_1116_nl;
  wire while_and_1117_nl;
  wire while_or_257_nl;
  wire while_and_1120_nl;
  wire while_and_1121_nl;
  wire PECore_PushAxiRsp_mux_24_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_nl;
  wire weight_mem_banks_load_store_1_for_else_else_or_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_4_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_6_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_8_nl;
  wire[7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_35_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_89_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_81_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_2_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl;
  wire mux_175_nl;
  wire nor_419_nl;
  wire nor_420_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_217_nl;
  wire mux_216_nl;
  wire mux_215_nl;
  wire or_581_nl;
  wire or_576_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_287_nl;
  wire mux_286_nl;
  wire mux_285_nl;
  wire or_665_nl;
  wire or_660_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_32_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl;
  wire nor_421_nl;
  wire mux_304_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl;
  wire PECore_UpdateFSM_switch_lp_mux1h_14_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl;
  wire PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl;
  wire PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_583_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_584_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_585_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_586_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_587_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_588_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_589_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_590_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_591_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_592_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_593_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_594_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_595_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_596_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_597_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_598_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_599_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_600_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_607_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_608_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_609_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_610_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_611_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_612_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_626_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_629_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_630_nl;
  wire mux_43_nl;
  wire mux_42_nl;
  wire mux_41_nl;
  wire and_699_nl;
  wire mux_59_nl;
  wire or_238_nl;
  wire or_234_nl;
  wire and_496_nl;
  wire and_495_nl;
  wire and_501_nl;
  wire and_500_nl;
  wire mux_106_nl;
  wire nor_320_nl;
  wire mux_108_nl;
  wire nor_321_nl;
  wire and_719_nl;
  wire nor_322_nl;
  wire or_374_nl;
  wire or_373_nl;
  wire and_722_nl;
  wire nor_323_nl;
  wire or_390_nl;
  wire or_389_nl;
  wire while_mux_1298_nl;
  wire or_495_nl;
  wire mux_159_nl;
  wire mux_158_nl;
  wire mux_157_nl;
  wire nand_8_nl;
  wire mux_156_nl;
  wire mux_155_nl;
  wire mux_154_nl;
  wire nand_7_nl;
  wire nor_358_nl;
  wire mux_166_nl;
  wire mux_165_nl;
  wire mux_164_nl;
  wire or_506_nl;
  wire or_505_nl;
  wire or_504_nl;
  wire nor_359_nl;
  wire mux_163_nl;
  wire mux_162_nl;
  wire mux_161_nl;
  wire or_499_nl;
  wire or_498_nl;
  wire mux_174_nl;
  wire mux_173_nl;
  wire mux_172_nl;
  wire mux_171_nl;
  wire nor_360_nl;
  wire nor_361_nl;
  wire nor_362_nl;
  wire nor_363_nl;
  wire mux_170_nl;
  wire mux_169_nl;
  wire mux_168_nl;
  wire nor_364_nl;
  wire nor_365_nl;
  wire nor_366_nl;
  wire nor_367_nl;
  wire mux_177_nl;
  wire mux_176_nl;
  wire or_534_nl;
  wire or_532_nl;
  wire nand_10_nl;
  wire nand_9_nl;
  wire mux_192_nl;
  wire mux_191_nl;
  wire mux_190_nl;
  wire mux_189_nl;
  wire mux_188_nl;
  wire mux_187_nl;
  wire mux_186_nl;
  wire mux_185_nl;
  wire mux_184_nl;
  wire mux_183_nl;
  wire mux_182_nl;
  wire mux_180_nl;
  wire mux_196_nl;
  wire mux_195_nl;
  wire mux_194_nl;
  wire or_545_nl;
  wire or_544_nl;
  wire or_543_nl;
  wire mux_200_nl;
  wire mux_199_nl;
  wire mux_198_nl;
  wire or_552_nl;
  wire or_551_nl;
  wire mux_206_nl;
  wire mux_205_nl;
  wire mux_204_nl;
  wire or_559_nl;
  wire or_558_nl;
  wire mux_203_nl;
  wire mux_202_nl;
  wire or_557_nl;
  wire or_556_nl;
  wire mux_201_nl;
  wire or_555_nl;
  wire or_548_nl;
  wire mux_214_nl;
  wire mux_213_nl;
  wire mux_212_nl;
  wire mux_211_nl;
  wire nor_368_nl;
  wire nor_369_nl;
  wire nor_370_nl;
  wire nor_371_nl;
  wire mux_210_nl;
  wire mux_209_nl;
  wire mux_208_nl;
  wire nor_372_nl;
  wire nor_373_nl;
  wire nor_374_nl;
  wire nor_375_nl;
  wire mux_219_nl;
  wire mux_218_nl;
  wire or_585_nl;
  wire or_583_nl;
  wire nand_12_nl;
  wire nand_11_nl;
  wire and_799_nl;
  wire mux_234_nl;
  wire mux_233_nl;
  wire mux_232_nl;
  wire mux_231_nl;
  wire mux_230_nl;
  wire mux_229_nl;
  wire mux_228_nl;
  wire mux_227_nl;
  wire mux_226_nl;
  wire mux_225_nl;
  wire mux_224_nl;
  wire or_589_nl;
  wire mux_222_nl;
  wire or_586_nl;
  wire or_603_nl;
  wire or_597_nl;
  wire mux_238_nl;
  wire mux_243_nl;
  wire mux_242_nl;
  wire or_607_nl;
  wire mux_241_nl;
  wire or_701_nl;
  wire or_606_nl;
  wire or_605_nl;
  wire mux_240_nl;
  wire or_702_nl;
  wire or_604_nl;
  wire mux_251_nl;
  wire mux_250_nl;
  wire mux_249_nl;
  wire mux_248_nl;
  wire or_614_nl;
  wire or_613_nl;
  wire or_612_nl;
  wire or_611_nl;
  wire mux_247_nl;
  wire mux_246_nl;
  wire mux_245_nl;
  wire or_610_nl;
  wire or_609_nl;
  wire or_608_nl;
  wire while_mux_1277_nl;
  wire mux_254_nl;
  wire mux_253_nl;
  wire or_621_nl;
  wire or_619_nl;
  wire mux_257_nl;
  wire mux_256_nl;
  wire nand_15_nl;
  wire mux_260_nl;
  wire mux_259_nl;
  wire nand_16_nl;
  wire mux_263_nl;
  wire mux_262_nl;
  wire or_623_nl;
  wire or_622_nl;
  wire mux_267_nl;
  wire mux_266_nl;
  wire mux_265_nl;
  wire or_628_nl;
  wire or_627_nl;
  wire or_626_nl;
  wire mux_270_nl;
  wire mux_269_nl;
  wire mux_268_nl;
  wire or_636_nl;
  wire or_635_nl;
  wire or_634_nl;
  wire mux_276_nl;
  wire mux_275_nl;
  wire mux_274_nl;
  wire or_643_nl;
  wire or_642_nl;
  wire mux_273_nl;
  wire mux_272_nl;
  wire or_641_nl;
  wire or_640_nl;
  wire mux_271_nl;
  wire or_639_nl;
  wire or_631_nl;
  wire mux_284_nl;
  wire mux_283_nl;
  wire mux_282_nl;
  wire mux_281_nl;
  wire nor_379_nl;
  wire nor_380_nl;
  wire nor_381_nl;
  wire nor_382_nl;
  wire mux_280_nl;
  wire mux_279_nl;
  wire mux_278_nl;
  wire nor_383_nl;
  wire nor_384_nl;
  wire nor_385_nl;
  wire nor_386_nl;
  wire mux_289_nl;
  wire mux_288_nl;
  wire or_669_nl;
  wire or_667_nl;
  wire while_mux_1255_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_625_nl;
  wire while_mux_1253_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_627_nl;
  wire mux_291_nl;
  wire mux_292_nl;
  wire mux_294_nl;
  wire mux_293_nl;
  wire or_680_nl;
  wire or_675_nl;
  wire or_690_nl;
  wire or_685_nl;
  wire mux_302_nl;
  wire mux_301_nl;
  wire mux_300_nl;
  wire mux_299_nl;
  wire or_703_nl;
  wire or_692_nl;
  wire mux_298_nl;
  wire or_704_nl;
  wire or_691_nl;
  wire mux_303_nl;
  wire weight_port_read_out_data_mux_48_nl;
  wire[6:0] weight_port_read_out_data_mux_75_nl;
  wire weight_port_read_out_data_mux_47_nl;
  wire[2:0] weight_port_read_out_data_mux_76_nl;
  wire[3:0] weight_port_read_out_data_mux_77_nl;
  wire weight_port_read_out_data_mux_46_nl;
  wire weight_port_read_out_data_mux_78_nl;
  wire[5:0] weight_port_read_out_data_mux_79_nl;
  wire[3:0] weight_port_read_out_data_mux_45_nl;
  wire[3:0] weight_port_read_out_data_mux_80_nl;
  wire weight_port_read_out_data_mux_44_nl;
  wire weight_port_read_out_data_mux_81_nl;
  wire[5:0] weight_port_read_out_data_mux_82_nl;
  wire weight_port_read_out_data_mux_43_nl;
  wire[6:0] weight_port_read_out_data_mux_83_nl;
  wire and_527_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl;
  wire weight_mem_banks_write_if_for_if_and_35_nl;
  wire weight_mem_banks_write_if_for_if_and_36_nl;
  wire weight_mem_banks_write_if_for_if_and_37_nl;
  wire weight_mem_banks_write_if_for_if_and_38_nl;
  wire weight_mem_banks_write_if_for_if_and_39_nl;
  wire weight_mem_banks_write_if_for_if_and_40_nl;
  wire weight_mem_banks_write_if_for_if_and_41_nl;
  wire weight_mem_banks_write_if_for_if_mux_7_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl;
  wire mux_151_nl;
  wire nor_412_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl;
  wire weight_mem_banks_write_if_for_if_and_28_nl;
  wire weight_mem_banks_write_if_for_if_and_29_nl;
  wire weight_mem_banks_write_if_for_if_and_30_nl;
  wire weight_mem_banks_write_if_for_if_and_31_nl;
  wire weight_mem_banks_write_if_for_if_and_32_nl;
  wire weight_mem_banks_write_if_for_if_and_33_nl;
  wire weight_mem_banks_write_if_for_if_and_34_nl;
  wire weight_mem_banks_write_if_for_if_mux_6_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl;
  wire mux_150_nl;
  wire nor_411_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl;
  wire weight_mem_banks_write_if_for_if_and_21_nl;
  wire weight_mem_banks_write_if_for_if_and_22_nl;
  wire weight_mem_banks_write_if_for_if_and_23_nl;
  wire weight_mem_banks_write_if_for_if_and_24_nl;
  wire weight_mem_banks_write_if_for_if_and_25_nl;
  wire weight_mem_banks_write_if_for_if_and_26_nl;
  wire weight_mem_banks_write_if_for_if_and_27_nl;
  wire weight_mem_banks_write_if_for_if_mux_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl;
  wire mux_149_nl;
  wire nor_410_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl;
  wire weight_mem_banks_write_if_for_if_and_14_nl;
  wire weight_mem_banks_write_if_for_if_and_15_nl;
  wire weight_mem_banks_write_if_for_if_and_16_nl;
  wire weight_mem_banks_write_if_for_if_and_17_nl;
  wire weight_mem_banks_write_if_for_if_and_18_nl;
  wire weight_mem_banks_write_if_for_if_and_19_nl;
  wire weight_mem_banks_write_if_for_if_and_20_nl;
  wire weight_mem_banks_write_if_for_if_mux_4_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl;
  wire mux_148_nl;
  wire nor_409_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl;
  wire weight_mem_banks_write_if_for_if_and_7_nl;
  wire weight_mem_banks_write_if_for_if_and_8_nl;
  wire weight_mem_banks_write_if_for_if_and_9_nl;
  wire weight_mem_banks_write_if_for_if_and_10_nl;
  wire weight_mem_banks_write_if_for_if_and_11_nl;
  wire weight_mem_banks_write_if_for_if_and_12_nl;
  wire weight_mem_banks_write_if_for_if_and_13_nl;
  wire weight_mem_banks_write_if_for_if_mux_3_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl;
  wire mux_147_nl;
  wire or_710_nl;
  wire mux_146_nl;
  wire or_406_nl;
  wire or_405_nl;
  wire nor_408_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl;
  wire weight_mem_banks_write_if_for_if_and_nl;
  wire weight_mem_banks_write_if_for_if_and_1_nl;
  wire weight_mem_banks_write_if_for_if_and_2_nl;
  wire weight_mem_banks_write_if_for_if_and_3_nl;
  wire weight_mem_banks_write_if_for_if_and_4_nl;
  wire weight_mem_banks_write_if_for_if_and_5_nl;
  wire weight_mem_banks_write_if_for_if_and_6_nl;
  wire weight_mem_banks_write_if_for_if_mux_2_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl;
  wire mux_145_nl;
  wire nor_406_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_1_nl;
  wire weight_mem_banks_write_if_for_if_mux_54_nl;
  wire mux_144_nl;
  wire nor_405_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_nl;
  wire weight_mem_banks_write_if_for_if_mux_53_nl;
  wire mux_143_nl;
  wire nor_404_nl;
  wire rva_out_reg_data_mux_20_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl;
  wire rva_out_reg_data_mux_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_22_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_18_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl;
  wire[5:0] PECore_DecodeAxiRead_switch_lp_mux_26_nl;
  wire rva_out_reg_data_mux_22_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_23_nl;
  wire PECore_PushAxiRsp_if_else_mux_17_nl;
  wire rva_out_reg_data_mux_24_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_24_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_20_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_27_nl;
  wire PECore_PushAxiRsp_if_else_mux_18_nl;
  wire rva_out_reg_data_mux_23_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl;
  wire mux_4_nl;
  wire mux_3_nl;
  wire mux_2_nl;
  wire or_5_nl;
  wire mux_58_nl;
  wire mux_61_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_8_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_38_nl;
  wire not_2208_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_15_nl;
  wire not_2209_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_39_nl;
  wire not_2210_nl;
  wire mux_69_nl;
  wire or_241_nl;
  wire[1:0] weight_mem_banks_load_store_for_else_mux1h_22_nl;
  wire not_2211_nl;
  wire[5:0] weight_mem_banks_load_store_for_else_mux1h_40_nl;
  wire not_2212_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_27_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_41_nl;
  wire not_2214_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_32_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_42_nl;
  wire not_2216_nl;
  wire mux1h_nl;
  wire[6:0] mux1h_8_nl;
  wire not_2301_nl;
  wire mux1h_2_nl;
  wire[6:0] mux1h_9_nl;
  wire not_2302_nl;
  wire mux1h_3_nl;
  wire mux1h_10_nl;
  wire[5:0] mux1h_11_nl;
  wire not_2303_nl;
  wire mux1h_4_nl;
  wire[2:0] mux1h_12_nl;
  wire not_2305_nl;
  wire[3:0] mux1h_13_nl;
  wire not_2306_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_136_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_137_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_64_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_87_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_65_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_80_nl;
  wire mux1h_5_nl;
  wire[6:0] mux1h_14_nl;
  wire not_2307_nl;
  wire[3:0] mux1h_6_nl;
  wire not_2308_nl;
  wire[3:0] mux1h_15_nl;
  wire not_2230_nl;
  wire mux1h_7_nl;
  wire mux1h_16_nl;
  wire[5:0] mux1h_17_nl;
  wire not_2309_nl;
  wire mux_1_nl;
  wire mux_886_nl;
  wire mux_885_nl;
  wire or_2319_nl;
  wire or_2318_nl;
  wire or_2317_nl;
  wire mux_887_nl;
  wire and_2185_nl;
  wire mux_890_nl;
  wire and_2186_nl;
  wire or_2327_nl;
  wire mux_895_nl;
  wire mux_894_nl;
  wire or_2340_nl;
  wire or_2339_nl;
  wire or_2338_nl;
  wire mux_896_nl;
  wire and_2188_nl;
  wire or_2341_nl;
  wire mux_899_nl;
  wire and_2189_nl;
  wire mux_902_nl;
  wire or_2355_nl;
  wire mux_905_nl;
  wire mux_908_nl;
  wire or_2371_nl;
  wire or_2369_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_19_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_25_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_30_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_28_nl;
  wire[3:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31_nl;
  wire[3:0] PECore_DecodeAxiRead_switch_lp_mux_29_nl;
  wire mux_742_nl;
  wire and_2070_nl;
  wire and_2071_nl;
  wire mux_780_nl;
  wire and_2095_nl;
  wire nor_1315_nl;
  wire mux_406_nl;
  wire nor_801_nl;
  wire nor_802_nl;
  wire mux_740_nl;
  wire and_2068_nl;
  wire nor_1261_nl;
  wire mux_408_nl;
  wire and_1895_nl;
  wire nor_805_nl;
  wire mux_862_nl;
  wire and_2165_nl;
  wire and_2166_nl;
  wire mux_806_nl;
  wire and_2113_nl;
  wire and_2114_nl;
  wire mux_590_nl;
  wire nor_1051_nl;
  wire nor_1052_nl;
  wire mux_540_nl;
  wire and_1953_nl;
  wire nor_983_nl;
  wire mux_390_nl;
  wire nor_779_nl;
  wire nor_780_nl;
  wire mux_418_nl;
  wire and_1900_nl;
  wire nor_818_nl;
  wire mux_508_nl;
  wire and_1939_nl;
  wire nor_941_nl;
  wire mux_456_nl;
  wire and_1914_nl;
  wire nor_869_nl;
  wire mux_628_nl;
  wire nor_1105_nl;
  wire nor_1106_nl;
  wire mux_674_nl;
  wire and_2028_nl;
  wire nor_1167_nl;
  wire mux_678_nl;
  wire and_2030_nl;
  wire nor_1173_nl;
  wire mux_850_nl;
  wire and_2152_nl;
  wire nor_1414_nl;
  wire mux_662_nl;
  wire nor_1149_nl;
  wire nor_1150_nl;
  wire mux_462_nl;
  wire nor_876_nl;
  wire nor_877_nl;
  wire mux_804_nl;
  wire and_2111_nl;
  wire nor_1350_nl;
  wire mux_544_nl;
  wire and_1954_nl;
  wire nor_988_nl;
  wire mux_530_nl;
  wire and_1948_nl;
  wire nor_969_nl;
  wire mux_526_nl;
  wire nor_963_nl;
  wire nor_964_nl;
  wire mux_846_nl;
  wire and_2148_nl;
  wire nor_1408_nl;
  wire mux_464_nl;
  wire nor_878_nl;
  wire nor_879_nl;
  wire mux_556_nl;
  wire and_1963_nl;
  wire nor_1006_nl;
  wire mux_610_nl;
  wire and_1995_nl;
  wire nor_1082_nl;
  wire mux_388_nl;
  wire and_1889_nl;
  wire nor_778_nl;
  wire mux_864_nl;
  wire and_2168_nl;
  wire and_2169_nl;
  wire mux_860_nl;
  wire and_2163_nl;
  wire nor_1427_nl;
  wire mux_856_nl;
  wire and_2158_nl;
  wire and_2159_nl;
  wire mux_554_nl;
  wire and_1962_nl;
  wire nor_1003_nl;
  wire mux_874_nl;
  wire and_2183_nl;
  wire and_2184_nl;
  wire mux_398_nl;
  wire nor_791_nl;
  wire nor_792_nl;
  wire mux_834_nl;
  wire and_2136_nl;
  wire nor_1392_nl;
  wire mux_792_nl;
  wire and_2101_nl;
  wire nor_1332_nl;
  wire mux_866_nl;
  wire and_2172_nl;
  wire nor_1434_nl;
  wire mux_826_nl;
  wire and_2130_nl;
  wire nor_1380_nl;
  wire mux_572_nl;
  wire and_1970_nl;
  wire nor_1027_nl;
  wire mux_648_nl;
  wire and_2015_nl;
  wire nor_1132_nl;
  wire mux_582_nl;
  wire and_1975_nl;
  wire nor_1041_nl;
  wire mux_436_nl;
  wire nor_842_nl;
  wire nor_843_nl;
  wire mux_380_nl;
  wire nor_765_nl;
  wire mux_379_nl;
  wire or_947_nl;
  wire or_945_nl;
  wire nor_766_nl;
  wire mux_402_nl;
  wire nor_797_nl;
  wire nor_798_nl;
  wire mux_726_nl;
  wire and_2057_nl;
  wire nor_1240_nl;
  wire mux_718_nl;
  wire nor_1227_nl;
  wire nor_1228_nl;
  wire mux_746_nl;
  wire and_2077_nl;
  wire nor_1268_nl;
  wire mux_372_nl;
  wire nor_754_nl;
  wire nor_755_nl;
  wire mux_772_nl;
  wire and_2089_nl;
  wire nor_1303_nl;
  wire mux_470_nl;
  wire nor_886_nl;
  wire nor_887_nl;
  wire mux_596_nl;
  wire and_1984_nl;
  wire nor_1061_nl;
  wire mux_642_nl;
  wire and_2013_nl;
  wire nor_1124_nl;
  wire mux_584_nl;
  wire and_1976_nl;
  wire nor_1044_nl;
  wire mux_636_nl;
  wire and_2011_nl;
  wire nor_1117_nl;
  wire mux_546_nl;
  wire and_1956_nl;
  wire nor_991_nl;
  wire mux_474_nl;
  wire and_1923_nl;
  wire nor_893_nl;
  wire mux_500_nl;
  wire nor_929_nl;
  wire nor_930_nl;
  wire mux_812_nl;
  wire and_2121_nl;
  wire nor_1360_nl;
  wire mux_810_nl;
  wire and_2120_nl;
  wire nor_1357_nl;
  wire mux_550_nl;
  wire and_1958_nl;
  wire nor_997_nl;
  wire mux_514_nl;
  wire and_1941_nl;
  wire nor_948_nl;
  wire mux_634_nl;
  wire and_2010_nl;
  wire nor_1114_nl;
  wire mux_664_nl;
  wire and_2022_nl;
  wire nor_1153_nl;
  wire mux_580_nl;
  wire and_1974_nl;
  wire nor_1038_nl;
  wire mux_702_nl;
  wire nor_1204_nl;
  wire nor_1205_nl;
  wire mux_468_nl;
  wire and_1920_nl;
  wire nor_885_nl;
  wire mux_844_nl;
  wire and_2147_nl;
  wire nor_1405_nl;
  wire mux_790_nl;
  wire and_2100_nl;
  wire nor_1329_nl;
  wire mux_606_nl;
  wire and_1991_nl;
  wire nor_1076_nl;
  wire mux_392_nl;
  wire and_1890_nl;
  wire nor_783_nl;
  wire mux_748_nl;
  wire and_2078_nl;
  wire nor_1271_nl;
  wire mux_752_nl;
  wire nor_1274_nl;
  wire nor_1275_nl;
  wire mux_708_nl;
  wire and_2046_nl;
  wire nor_1214_nl;
  wire mux_598_nl;
  wire and_1985_nl;
  wire nor_1064_nl;
  wire mux_758_nl;
  wire nor_1282_nl;
  wire nor_1283_nl;
  wire mux_506_nl;
  wire and_1938_nl;
  wire nor_938_nl;
  wire mux_426_nl;
  wire and_1904_nl;
  wire nor_829_nl;
  wire mux_446_nl;
  wire nor_855_nl;
  wire nor_856_nl;
  wire mux_680_nl;
  wire and_2031_nl;
  wire nor_1176_nl;
  wire mux_480_nl;
  wire and_1925_nl;
  wire nor_901_nl;
  wire mux_516_nl;
  wire and_1942_nl;
  wire nor_951_nl;
  wire mux_412_nl;
  wire and_1898_nl;
  wire nor_811_nl;
  wire mux_494_nl;
  wire nor_921_nl;
  wire nor_922_nl;
  wire mux_444_nl;
  wire and_1910_nl;
  wire nor_854_nl;
  wire mux_424_nl;
  wire and_1902_nl;
  wire nor_826_nl;
  wire mux_666_nl;
  wire and_2024_nl;
  wire nor_1156_nl;
  wire mux_452_nl;
  wire and_1913_nl;
  wire nor_864_nl;
  wire mux_578_nl;
  wire and_1973_nl;
  wire nor_1035_nl;
  wire mux_366_nl;
  wire nor_745_nl;
  wire nor_746_nl;
  wire mux_442_nl;
  wire and_1909_nl;
  wire nor_851_nl;
  wire mux_486_nl;
  wire and_1929_nl;
  wire nor_910_nl;
  wire mux_638_nl;
  wire nor_1118_nl;
  wire nor_1119_nl;
  wire mux_808_nl;
  wire and_2116_nl;
  wire and_2117_nl;
  wire mux_694_nl;
  wire nor_1193_nl;
  wire nor_1194_nl;
  wire mux_552_nl;
  wire and_1959_nl;
  wire nor_1000_nl;
  wire mux_872_nl;
  wire and_2180_nl;
  wire and_2181_nl;
  wire mux_778_nl;
  wire and_2094_nl;
  wire nor_1312_nl;
  wire mux_458_nl;
  wire and_1916_nl;
  wire nor_872_nl;
  wire mux_542_nl;
  wire nor_984_nl;
  wire nor_985_nl;
  wire mux_820_nl;
  wire and_2125_nl;
  wire nor_1371_nl;
  wire mux_832_nl;
  wire and_2133_nl;
  wire nor_1389_nl;
  wire mux_750_nl;
  wire nor_1272_nl;
  wire nor_1273_nl;
  wire mux_738_nl;
  wire and_2067_nl;
  wire nor_1258_nl;
  wire mux_454_nl;
  wire nor_865_nl;
  wire nor_866_nl;
  wire mux_588_nl;
  wire and_1980_nl;
  wire nor_1050_nl;
  wire mux_386_nl;
  wire nor_774_nl;
  wire nor_775_nl;
  wire mux_496_nl;
  wire nor_924_nl;
  wire nor_925_nl;
  wire mux_394_nl;
  wire and_1892_nl;
  wire nor_786_nl;
  wire mux_732_nl;
  wire and_2062_nl;
  wire nor_1249_nl;
  wire mux_570_nl;
  wire and_1969_nl;
  wire nor_1024_nl;
  wire mux_612_nl;
  wire and_1996_nl;
  wire nor_1085_nl;
  wire mux_728_nl;
  wire and_2058_nl;
  wire nor_1243_nl;
  wire mux_858_nl;
  wire and_2162_nl;
  wire nor_1424_nl;
  wire mux_532_nl;
  wire and_1949_nl;
  wire nor_972_nl;
  wire mux_698_nl;
  wire and_2041_nl;
  wire nor_1200_nl;
  wire mux_660_nl;
  wire and_2021_nl;
  wire nor_1148_nl;
  wire mux_818_nl;
  wire and_2124_nl;
  wire nor_1368_nl;
  wire mux_828_nl;
  wire and_2131_nl;
  wire nor_1383_nl;
  wire mux_736_nl;
  wire and_2064_nl;
  wire nor_1255_nl;
  wire mux_870_nl;
  wire and_2177_nl;
  wire and_2178_nl;
  wire mux_574_nl;
  wire nor_1028_nl;
  wire nor_1029_nl;
  wire mux_566_nl;
  wire nor_1017_nl;
  wire nor_1018_nl;
  wire mux_378_nl;
  wire nor_763_nl;
  wire nor_764_nl;
  wire mux_374_nl;
  wire nor_757_nl;
  wire nor_758_nl;
  wire mux_766_nl;
  wire nor_1293_nl;
  wire nor_1294_nl;
  wire mux_836_nl;
  wire and_2137_nl;
  wire nor_1395_nl;
  wire mux_754_nl;
  wire and_2080_nl;
  wire nor_1278_nl;
  wire mux_488_nl;
  wire and_1930_nl;
  wire nor_913_nl;
  wire mux_548_nl;
  wire and_1957_nl;
  wire nor_994_nl;
  wire mux_400_nl;
  wire nor_794_nl;
  wire nor_795_nl;
  wire mux_434_nl;
  wire nor_840_nl;
  wire nor_841_nl;
  wire mux_784_nl;
  wire and_2096_nl;
  wire nor_1320_nl;
  wire mux_576_nl;
  wire and_1971_nl;
  wire nor_1032_nl;
  wire mux_504_nl;
  wire and_1936_nl;
  wire nor_935_nl;
  wire mux_616_nl;
  wire and_2001_nl;
  wire and_2002_nl;
  wire mux_370_nl;
  wire nor_751_nl;
  wire nor_752_nl;
  wire mux_558_nl;
  wire nor_1007_nl;
  wire nor_1008_nl;
  wire mux_868_nl;
  wire and_2174_nl;
  wire and_2175_nl;
  wire mux_518_nl;
  wire nor_952_nl;
  wire nor_953_nl;
  wire mux_478_nl;
  wire nor_897_nl;
  wire nor_898_nl;
  wire mux_798_nl;
  wire and_2106_nl;
  wire nor_1341_nl;
  wire mux_690_nl;
  wire and_2037_nl;
  wire nor_1189_nl;
  wire mux_396_nl;
  wire and_1893_nl;
  wire nor_789_nl;
  wire mux_448_nl;
  wire nor_857_nl;
  wire nor_858_nl;
  wire mux_802_nl;
  wire and_2110_nl;
  wire nor_1347_nl;
  wire mux_814_nl;
  wire nor_1361_nl;
  wire nor_1362_nl;
  wire mux_604_nl;
  wire and_1990_nl;
  wire nor_1073_nl;
  wire mux_490_nl;
  wire and_1933_nl;
  wire nor_916_nl;
  wire mux_822_nl;
  wire and_2126_nl;
  wire nor_1374_nl;
  wire mux_716_nl;
  wire and_2052_nl;
  wire nor_1226_nl;
  wire mux_472_nl;
  wire and_1921_nl;
  wire nor_890_nl;
  wire mux_512_nl;
  wire nor_944_nl;
  wire nor_945_nl;
  wire mux_524_nl;
  wire and_1946_nl;
  wire nor_962_nl;
  wire mux_520_nl;
  wire and_1943_nl;
  wire nor_956_nl;
  wire mux_644_nl;
  wire and_2014_nl;
  wire nor_1127_nl;
  wire mux_670_nl;
  wire nor_1160_nl;
  wire nor_1161_nl;
  wire mux_712_nl;
  wire and_2048_nl;
  wire nor_1220_nl;
  wire mux_676_nl;
  wire and_2029_nl;
  wire nor_1170_nl;
  wire mux_768_nl;
  wire and_2086_nl;
  wire nor_1297_nl;
  wire mux_840_nl;
  wire and_2142_nl;
  wire and_2143_nl;
  wire mux_498_nl;
  wire nor_927_nl;
  wire nor_928_nl;
  wire mux_538_nl;
  wire and_1952_nl;
  wire nor_980_nl;
  wire mux_658_nl;
  wire and_2020_nl;
  wire nor_1145_nl;
  wire mux_704_nl;
  wire and_2043_nl;
  wire nor_1208_nl;
  wire mux_368_nl;
  wire nor_748_nl;
  wire nor_749_nl;
  wire mux_422_nl;
  wire nor_822_nl;
  wire nor_823_nl;
  wire mux_730_nl;
  wire and_2061_nl;
  wire nor_1246_nl;
  wire mux_696_nl;
  wire and_2039_nl;
  wire nor_1197_nl;
  wire mux_430_nl;
  wire nor_834_nl;
  wire nor_835_nl;
  wire mux_632_nl;
  wire and_2008_nl;
  wire nor_1111_nl;
  wire mux_688_nl;
  wire nor_1185_nl;
  wire nor_1186_nl;
  wire mux_682_nl;
  wire and_2034_nl;
  wire nor_1179_nl;
  wire mux_466_nl;
  wire and_1919_nl;
  wire nor_882_nl;
  wire mux_668_nl;
  wire and_2025_nl;
  wire nor_1159_nl;
  wire mux_710_nl;
  wire and_2047_nl;
  wire nor_1217_nl;
  wire mux_722_nl;
  wire and_2055_nl;
  wire nor_1234_nl;
  wire mux_724_nl;
  wire and_2056_nl;
  wire nor_1237_nl;
  wire mux_652_nl;
  wire and_2018_nl;
  wire nor_1138_nl;
  wire mux_782_nl;
  wire nor_1316_nl;
  wire nor_1317_nl;
  wire mux_460_nl;
  wire and_1917_nl;
  wire nor_875_nl;
  wire mux_684_nl;
  wire and_2035_nl;
  wire nor_1182_nl;
  wire mux_770_nl;
  wire and_2088_nl;
  wire nor_1300_nl;
  wire mux_404_nl;
  wire nor_799_nl;
  wire nor_800_nl;
  wire mux_450_nl;
  wire and_1912_nl;
  wire nor_861_nl;
  wire mux_838_nl;
  wire and_2139_nl;
  wire and_2140_nl;
  wire mux_568_nl;
  wire and_1967_nl;
  wire nor_1021_nl;
  wire mux_586_nl;
  wire and_1979_nl;
  wire nor_1047_nl;
  wire mux_622_nl;
  wire nor_1097_nl;
  wire nor_1098_nl;
  wire mux_564_nl;
  wire and_1966_nl;
  wire nor_1016_nl;
  wire mux_384_nl;
  wire nor_771_nl;
  wire nor_772_nl;
  wire mux_654_nl;
  wire nor_1139_nl;
  wire nor_1140_nl;
  wire mux_842_nl;
  wire and_2146_nl;
  wire nor_1402_nl;
  wire mux_756_nl;
  wire and_2081_nl;
  wire nor_1281_nl;
  wire mux_476_nl;
  wire and_1924_nl;
  wire nor_896_nl;
  wire mux_672_nl;
  wire and_2026_nl;
  wire nor_1164_nl;
  wire mux_646_nl;
  wire nor_1128_nl;
  wire nor_1129_nl;
  wire mux_854_nl;
  wire and_2155_nl;
  wire and_2156_nl;
  wire mux_620_nl;
  wire and_2006_nl;
  wire nor_1095_nl;
  wire mux_692_nl;
  wire and_2038_nl;
  wire nor_1192_nl;
  wire mux_714_nl;
  wire and_2051_nl;
  wire nor_1223_nl;
  wire mux_502_nl;
  wire nor_931_nl;
  wire nor_932_nl;
  wire mux_376_nl;
  wire nor_760_nl;
  wire nor_761_nl;
  wire mux_614_nl;
  wire and_1998_nl;
  wire and_1999_nl;
  wire mux_618_nl;
  wire and_2005_nl;
  wire nor_1092_nl;
  wire mux_528_nl;
  wire nor_965_nl;
  wire nor_966_nl;
  wire mux_414_nl;
  wire nor_812_nl;
  wire nor_813_nl;
  wire mux_816_nl;
  wire and_2122_nl;
  wire nor_1365_nl;
  wire mux_640_nl;
  wire nor_1120_nl;
  wire nor_1121_nl;
  wire mux_630_nl;
  wire nor_1107_nl;
  wire nor_1108_nl;
  wire mux_438_nl;
  wire nor_844_nl;
  wire nor_845_nl;
  wire mux_848_nl;
  wire and_2149_nl;
  wire nor_1411_nl;
  wire mux_706_nl;
  wire and_2045_nl;
  wire nor_1211_nl;
  wire mux_796_nl;
  wire and_2105_nl;
  wire nor_1338_nl;
  wire mux_776_nl;
  wire and_2091_nl;
  wire nor_1309_nl;
  wire mux_382_nl;
  wire nor_768_nl;
  wire nor_769_nl;
  wire mux_428_nl;
  wire and_1905_nl;
  wire nor_832_nl;
  wire mux_536_nl;
  wire and_1950_nl;
  wire nor_977_nl;
  wire mux_608_nl;
  wire and_1992_nl;
  wire nor_1079_nl;
  wire mux_416_nl;
  wire nor_814_nl;
  wire nor_815_nl;
  wire mux_744_nl;
  wire and_2073_nl;
  wire and_2074_nl;
  wire mux_762_nl;
  wire and_2084_nl;
  wire nor_1289_nl;
  wire mux_510_nl;
  wire nor_942_nl;
  wire nor_943_nl;
  wire mux_522_nl;
  wire and_1945_nl;
  wire nor_959_nl;
  wire mux_592_nl;
  wire and_1981_nl;
  wire nor_1055_nl;
  wire mux_626_nl;
  wire nor_1103_nl;
  wire nor_1104_nl;
  wire mux_760_nl;
  wire and_2082_nl;
  wire nor_1286_nl;
  wire mux_560_nl;
  wire nor_1009_nl;
  wire nor_1010_nl;
  wire mux_700_nl;
  wire and_2042_nl;
  wire nor_1203_nl;
  wire mux_656_nl;
  wire nor_1141_nl;
  wire nor_1142_nl;
  wire mux_786_nl;
  wire and_2098_nl;
  wire nor_1323_nl;
  wire mux_830_nl;
  wire and_2132_nl;
  wire nor_1386_nl;
  wire mux_594_nl;
  wire and_1983_nl;
  wire nor_1058_nl;
  wire mux_794_nl;
  wire and_2104_nl;
  wire nor_1335_nl;
  wire mux_788_nl;
  wire and_2099_nl;
  wire nor_1326_nl;
  wire mux_764_nl;
  wire and_2085_nl;
  wire nor_1292_nl;
  wire mux_650_nl;
  wire and_2017_nl;
  wire nor_1135_nl;
  wire mux_734_nl;
  wire and_2063_nl;
  wire nor_1252_nl;
  wire mux_410_nl;
  wire and_1897_nl;
  wire nor_808_nl;
  wire mux_774_nl;
  wire and_2090_nl;
  wire nor_1306_nl;
  wire mux_562_nl;
  wire and_1965_nl;
  wire nor_1013_nl;
  wire mux_440_nl;
  wire and_1907_nl;
  wire nor_848_nl;
  wire mux_824_nl;
  wire and_2127_nl;
  wire nor_1377_nl;
  wire mux_800_nl;
  wire and_2107_nl;
  wire nor_1344_nl;
  wire mux_852_nl;
  wire and_2153_nl;
  wire nor_1417_nl;
  wire mux_686_nl;
  wire nor_1183_nl;
  wire nor_1184_nl;
  wire mux_484_nl;
  wire and_1928_nl;
  wire nor_907_nl;
  wire mux_624_nl;
  wire nor_1100_nl;
  wire nor_1101_nl;
  wire mux_720_nl;
  wire and_2053_nl;
  wire nor_1231_nl;
  wire mux_602_nl;
  wire and_1989_nl;
  wire nor_1070_nl;
  wire mux_600_nl;
  wire and_1986_nl;
  wire nor_1067_nl;
  wire mux_432_nl;
  wire nor_837_nl;
  wire nor_838_nl;
  wire mux_420_nl;
  wire and_1901_nl;
  wire nor_821_nl;
  wire mux_534_nl;
  wire nor_973_nl;
  wire nor_974_nl;
  wire mux_492_nl;
  wire and_1934_nl;
  wire nor_919_nl;
  wire mux_482_nl;
  wire and_1927_nl;
  wire nor_904_nl;
  wire mux_364_nl;
  wire nor_742_nl;
  wire mux_363_nl;
  wire or_900_nl;
  wire or_899_nl;
  wire nor_743_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (~ reg_rva_in_reg_rw_sva_2_cse);
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0];
  wire  nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a = PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2
      & reg_rva_in_reg_rw_sva_2_cse;
  wire [2:0] nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s = weight_write_addrs_lpi_1_dfm_1_2[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s = {(weight_read_addrs_6_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_4[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s = weight_read_addrs_7_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s = {(weight_read_addrs_2_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s = {(weight_read_addrs_4_14_2_lpi_1_dfm_1_1[0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[1:0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s = weight_read_addrs_3_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s = weight_read_addrs_5_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s = weight_read_addrs_1_lpi_1_dfm_1_1[2:0];
  wire [255:0] nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff;
  assign nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff
      = {16'b0000000000000000 , act_port_reg_data_239_224_sva_dfm_1_2 , 16'b0000000000000000
      , act_port_reg_data_207_192_sva_dfm_1_2 , 16'b0000000000000000 , act_port_reg_data_175_160_sva_dfm_1_2
      , 16'b0000000000000000 , act_port_reg_data_143_128_sva_dfm_1_2 , 16'b0000000000000000
      , act_port_reg_data_111_96_sva_dfm_1_2 , 16'b0000000000000000 , act_port_reg_data_79_64_sva_dfm_1_1
      , 16'b0000000000000000 , act_port_reg_data_47_32_sva_dfm_1_2 , 16'b0000000000000000
      , act_port_reg_data_15_0_sva_dfm_1_2};
  wire weight_port_read_out_data_mux_4_nl;
  wire weight_port_read_out_data_mux_86_nl;
  wire weight_port_read_out_data_mux_2_nl;
  wire weight_port_read_out_data_mux_85_nl;
  wire weight_port_read_out_data_mux_nl;
  wire weight_port_read_out_data_mux_84_nl;
  wire [63:0] nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign weight_port_read_out_data_mux_86_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_16_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign weight_port_read_out_data_mux_4_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2,
      weight_port_read_out_data_mux_86_nl, fsm_output);
  assign weight_port_read_out_data_mux_85_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_15_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign weight_port_read_out_data_mux_2_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2,
      weight_port_read_out_data_mux_85_nl, fsm_output);
  assign weight_port_read_out_data_mux_84_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_14_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign weight_port_read_out_data_mux_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2,
      weight_port_read_out_data_mux_84_nl, fsm_output);
  assign nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun
      = {rva_out_reg_data_63_sva_dfm_4_5 , rva_out_reg_data_62_56_sva_dfm_4_5 , rva_out_reg_data_55_48_sva_dfm_4_5_7_4
      , rva_out_reg_data_55_48_sva_dfm_4_5_3_0 , rva_out_reg_data_47_sva_dfm_4_5
      , rva_out_reg_data_46_40_sva_dfm_4_5_6_4 , rva_out_reg_data_46_40_sva_dfm_4_5_3_0
      , rva_out_reg_data_39_36_sva_dfm_4_5_3 , rva_out_reg_data_39_36_sva_dfm_4_5_2
      , rva_out_reg_data_39_36_sva_dfm_4_5_1_0 , rva_out_reg_data_35_32_sva_dfm_4_5
      , PECore_PushAxiRsp_if_mux1h_17 , PECore_PushAxiRsp_if_mux1h_16_5_3 , PECore_PushAxiRsp_if_mux1h_16_2_0
      , PECore_PushAxiRsp_if_mux1h_15 , PECore_PushAxiRsp_if_mux1h_14_6 , PECore_PushAxiRsp_if_mux1h_14_5
      , PECore_PushAxiRsp_if_mux1h_14_4 , PECore_PushAxiRsp_if_mux1h_14_3_0 , weight_port_read_out_data_mux_4_nl
      , PECore_PushAxiRsp_if_mux1h_12_6 , PECore_PushAxiRsp_if_mux1h_12_5_0 , weight_port_read_out_data_mux_2_nl
      , PECore_PushAxiRsp_if_mux1h_10_6 , PECore_PushAxiRsp_if_mux1h_10_5_0 , weight_port_read_out_data_mux_nl};
  PECore_mgc_muladd1 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_cst(32'sd1),
  .signd_cst(32'sd0),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd11),
  .add_axb(32'sd1),
  .add_c(32'sd1),
  .add_d(32'sd1),
  .use_const(32'sd1)) PEManager_15U_GetWeightAddr_else_acc_4_cmp (
      .a(pe_config_output_counter_sva),
      .b(pe_manager_num_input_sva),
      .c(pe_config_input_counter_sva),
      .cst(1'b0),
      .z(PEManager_15U_GetWeightAddr_else_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_for_1_lshift_rg (
      .a(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a),
      .s(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_write_arbxbar_xbar_for_lshift_rg (
      .a(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a),
      .s(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s[2:0]),
      .z(weight_mem_write_arbxbar_xbar_for_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi PECore_PECoreRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(fsm_output)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi PECore_PECoreRun_input_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_oswt_pff(and_524_rmff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi PECore_PECoreRun_act_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(reg_act_port_Push_mioi_iswt0_cse),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff(nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun_pff[255:0]),
      .act_port_Push_mioi_oswt_pff(and_526_rmff)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi PECore_PECoreRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_oswt_pff(and_524_rmff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi PECore_PECoreRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun[63:0]),
      .rva_out_Push_mioi_oswt_pff(and_522_cse)
    );
  PECore_PECore_PECoreRun_wait_dp PECore_PECoreRun_wait_dp_inst (
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_en(Datapath_for_4_ProductSum_for_acc_5_cmp_21_en),
      .PECoreRun_wen(PECoreRun_wen),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg(and_520_rmff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg(and_517_rmff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg(and_514_rmff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg(and_511_rmff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg(and_508_rmff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg(and_505_rmff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg(and_502_rmff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg(and_497_rmff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_cgo(reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_31_cse),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg(and_489_rmff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_21(reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_21_cse),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_unreg_21(and_492_rmff)
    );
  PECore_PECore_PECoreRun_staller PECore_PECoreRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp)
    );
  PECore_PECore_PECoreRun_PECoreRun_fsm PECore_PECoreRun_PECoreRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .fsm_output(fsm_output)
    );
  assign weight_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_84);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign weight_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_84);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign weight_mem_banks_read_1_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_85);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign weight_mem_banks_read_1_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_85);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign weight_mem_banks_read_1_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_86);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 );
  assign weight_mem_banks_read_1_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_86);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign weight_mem_banks_read_1_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_87);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 );
  assign weight_mem_banks_read_1_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_87);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign weight_mem_banks_read_1_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_89);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 );
  assign weight_mem_banks_read_1_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_89);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign weight_mem_banks_read_1_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_90);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 );
  assign weight_mem_banks_read_1_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_90);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign weight_mem_banks_read_1_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_81);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 );
  assign weight_mem_banks_read_1_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_81);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign weight_mem_banks_read_1_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_83);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 );
  assign weight_mem_banks_read_1_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_83);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign weight_mem_banks_write_if_for_if_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_170);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 );
  assign weight_mem_banks_write_if_for_if_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_170);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign weight_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_171);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 );
  assign weight_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_171);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign weight_mem_banks_write_if_for_if_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_173);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 );
  assign weight_mem_banks_write_if_for_if_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_173);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1
      = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1
      = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign weight_mem_banks_read_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_174);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 );
  assign weight_mem_banks_read_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_174);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign weight_mem_banks_write_if_for_if_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_176);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 );
  assign weight_mem_banks_write_if_for_if_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_176);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2
      = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2
      = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign weight_mem_banks_read_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_177);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 );
  assign weight_mem_banks_read_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_177);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign weight_mem_banks_write_if_for_if_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_179);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 );
  assign weight_mem_banks_write_if_for_if_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_179);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3
      = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3
      = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign weight_mem_banks_read_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_180);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 );
  assign weight_mem_banks_read_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_180);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign weight_mem_banks_write_if_for_if_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_182);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 );
  assign weight_mem_banks_write_if_for_if_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_182);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4
      = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4
      = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign weight_mem_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_183);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 );
  assign weight_mem_banks_read_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_183);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign weight_mem_banks_write_if_for_if_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_185);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 );
  assign weight_mem_banks_write_if_for_if_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_185);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5
      = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5
      = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign weight_mem_banks_read_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_186);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 );
  assign weight_mem_banks_read_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_186);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign weight_mem_banks_write_if_for_if_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_187);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 );
  assign weight_mem_banks_write_if_for_if_mux_33_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_187);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6
      = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6
      = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign weight_mem_banks_read_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_188);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 );
  assign weight_mem_banks_read_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_188);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign weight_mem_banks_write_if_for_if_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_190);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 );
  assign weight_mem_banks_write_if_for_if_mux_37_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_190);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7
      = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7
      = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign weight_mem_banks_read_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_191);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 );
  assign weight_mem_banks_read_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_191);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign input_mem_banks_write_1_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_201);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 );
  assign input_mem_banks_write_1_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_201);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8
      = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_3 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8
      = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign input_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_198);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 );
  assign input_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_198);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign input_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_208);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 );
  assign input_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_208);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9
      = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_1 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9
      = input_mem_banks_write_if_for_if_mux_1_cse;
  assign input_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_211);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 );
  assign input_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_211);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign and_489_rmff = (and_dcpl_480 | (PECore_RunMac_PECore_RunMac_if_and_svs_st_5
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7) | and_dcpl_476) & fsm_output;
  assign and_492_rmff = (and_dcpl_480 | (while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_8) | and_dcpl_476) & fsm_output;
  assign or_705_nl = (while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
      & (~ weight_mem_run_3_for_5_and_132_itm_1)) | mux_tmp_99;
  assign nand_2_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~((~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3)
      | weight_mem_run_3_for_5_and_132_itm_1)) | mux_tmp_99)));
  assign mux_100_nl = MUX_s_1_2_2(mux_tmp_99, nand_2_nl, while_stage_0_7);
  assign mux_101_nl = MUX_s_1_2_2(or_705_nl, mux_100_nl, weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign and_497_rmff = (mux_101_nl | and_dcpl_486) & fsm_output;
  assign or_347_nl = (while_stage_0_7 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1)
      & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3)
      | mux_tmp_103;
  assign nand_4_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & (~((~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3)))
      | mux_tmp_103)));
  assign mux_104_nl = MUX_s_1_2_2(mux_tmp_103, nand_4_nl, while_stage_0_7);
  assign mux_105_nl = MUX_s_1_2_2(or_347_nl, mux_104_nl, weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign and_502_rmff = (mux_105_nl | and_dcpl_489) & fsm_output;
  assign or_353_nl = (weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      & while_stage_0_5) | not_tmp_264;
  assign or_351_nl = (((weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]) | weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1)
      & while_stage_0_5) | not_tmp_264;
  assign mux_107_nl = MUX_s_1_2_2(or_353_nl, or_351_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_505_rmff = (mux_107_nl | and_dcpl_185) & fsm_output;
  assign or_360_nl = (or_708_cse & while_stage_0_5) | not_tmp_267;
  assign or_357_nl = (((weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]) | weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1)
      & while_stage_0_5) | not_tmp_267;
  assign mux_109_nl = MUX_s_1_2_2(or_360_nl, or_357_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_508_rmff = (mux_109_nl | and_dcpl_182) & fsm_output;
  assign or_367_nl = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      | not_tmp_270;
  assign or_365_nl = (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]) | PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3
      | not_tmp_270;
  assign mux_111_nl = MUX_s_1_2_2(or_367_nl, or_365_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_112_nl = MUX_s_1_2_2(not_tmp_270, mux_111_nl, while_stage_0_5);
  assign and_511_rmff = (mux_112_nl | and_dcpl_179) & fsm_output;
  assign or_375_nl = (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]) | PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
  assign mux_116_nl = MUX_s_1_2_2(not_tmp_274, mux_tmp_113, or_375_nl);
  assign mux_117_nl = MUX_s_1_2_2(not_tmp_274, mux_116_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_370_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]) | PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
  assign mux_115_nl = MUX_s_1_2_2(not_tmp_274, mux_tmp_113, or_370_nl);
  assign mux_118_nl = MUX_s_1_2_2(mux_117_nl, mux_115_nl, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse);
  assign and_514_rmff = (mux_118_nl | and_dcpl_176) & fsm_output;
  assign or_383_nl = PECore_RunMac_PECore_RunMac_if_and_svs_st_3 | PECore_UpdateFSM_switch_lp_equal_tmp_2_3
      | not_tmp_277;
  assign mux_121_nl = MUX_s_1_2_2(not_tmp_277, or_383_nl, and_882_cse);
  assign or_381_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_3 | PECore_UpdateFSM_switch_lp_equal_tmp_2_3
      | not_tmp_277;
  assign mux_120_nl = MUX_s_1_2_2(not_tmp_277, or_381_nl, while_stage_0_5);
  assign mux_122_nl = MUX_s_1_2_2(mux_121_nl, mux_120_nl, weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse);
  assign and_517_rmff = (mux_122_nl | and_dcpl_173) & fsm_output;
  assign or_391_nl = PECore_RunFSM_switch_lp_equal_tmp_1_2 | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
  assign mux_126_nl = MUX_s_1_2_2(not_tmp_281, mux_tmp_123, or_391_nl);
  assign mux_127_nl = MUX_s_1_2_2(not_tmp_281, mux_126_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_386_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | PECore_RunFSM_switch_lp_equal_tmp_1_2 | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
  assign mux_125_nl = MUX_s_1_2_2(not_tmp_281, mux_tmp_123, or_386_nl);
  assign mux_128_nl = MUX_s_1_2_2(mux_127_nl, mux_125_nl, weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse);
  assign and_520_rmff = (mux_128_nl | and_dcpl_170) & fsm_output;
  assign and_990_itm = PECore_UpdateFSM_switch_lp_nor_7_itm_1 & PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      & pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign and_702_itm = pe_config_is_zero_first_sva & PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      & pe_manager_zero_active_sva;
  assign and_709_cse = PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign mux_924_nl = MUX_s_1_2_2(and_990_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_702_itm);
  assign and_708_nl = start_PopNB_mioi_data_rsc_z_mxwt & start_PopNB_mioi_return_rsc_z_mxwt
      & PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign mux_137_nl = MUX_s_1_2_2(mux_924_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_708_nl);
  assign mux_322_nl = MUX_s_1_2_2(and_990_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_702_itm);
  assign mux_133_nl = MUX_s_1_2_2(mux_322_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_709_cse);
  assign mux_138_nl = MUX_s_1_2_2(mux_137_nl, mux_133_nl, or_220_cse);
  assign mux_926_nl = MUX_s_1_2_2(and_990_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_702_itm);
  assign mux_925_nl = MUX_s_1_2_2(mux_926_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_709_cse);
  assign or_218_nl = pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]);
  assign mux_134_nl = MUX_s_1_2_2(mux_925_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_218_nl);
  assign or_217_nl = (state_2_1_sva!=2'b10) | state_0_sva;
  assign mux_135_nl = MUX_s_1_2_2(mux_134_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_217_nl);
  assign mux_136_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_nor_7_itm_1, mux_135_nl,
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign mux_139_nl = MUX_s_1_2_2(mux_138_nl, mux_136_nl, PECore_UpdateFSM_switch_lp_equal_tmp_5_1);
  assign mux_140_nl = MUX_s_1_2_2(mux_139_nl, state_0_sva, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_141_nl = MUX_s_1_2_2(or_220_cse, mux_140_nl, while_stage_0_3);
  assign or_216_nl = while_stage_0_3 | (state_2_1_sva!=2'b00) | state_0_sva;
  assign or_215_nl = (state_2_1_sva_dfm_1!=2'b00);
  assign mux_142_cse = MUX_s_1_2_2(mux_141_nl, or_216_nl, or_215_nl);
  assign and_524_rmff = (~ mux_142_cse) & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign and_526_rmff = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10)
      & while_stage_0_12 & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10;
  assign PECore_DecodeAxiRead_switch_lp_and_2_cse = PECoreRun_wen & and_dcpl_6;
  assign rva_out_reg_data_and_14_cse = PECoreRun_wen & and_dcpl_6 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_9) & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9));
  assign rva_out_reg_data_and_90_enex5 = rva_out_reg_data_and_14_cse & reg_rva_out_reg_data_30_25_sva_dfm_7_enexo;
  assign rva_out_reg_data_and_17_cse = PECoreRun_wen & and_dcpl_5;
  assign rva_out_reg_data_and_91_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_92_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo;
  assign input_mem_banks_read_read_data_and_cse = PECoreRun_wen & and_dcpl_5 & (~
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7) & input_read_req_valid_lpi_1_dfm_1_9;
  assign weight_port_read_out_data_and_64_cse = PECoreRun_wen & and_dcpl_4 & (~ rva_in_reg_rw_sva_st_1_9)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
  assign rva_out_reg_data_and_cse = PECoreRun_wen & (~((~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
      & while_stage_0_12)) | rva_in_reg_rw_sva_10 | (~ fsm_output)));
  assign input_mem_banks_read_read_data_and_31_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_32_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_33_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo;
  assign input_mem_banks_read_read_data_and_34_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo;
  assign rva_in_reg_rw_and_cse = PECoreRun_wen & while_stage_0_11;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_cse = PECoreRun_wen & and_dcpl_4
      & (~(rva_in_reg_rw_sva_st_1_9 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7))
      & (~(input_read_req_valid_lpi_1_dfm_1_9 | rva_in_reg_rw_sva_9)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
  assign act_port_reg_data_and_cse = PECoreRun_wen & and_dcpl_22 & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  assign act_port_reg_data_and_30_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_15_0_sva_dfm_1_1_enexo;
  assign act_port_reg_data_and_31_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_239_224_sva_dfm_1_1_enexo;
  assign act_port_reg_data_and_32_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_47_32_sva_dfm_1_1_enexo;
  assign act_port_reg_data_and_33_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_207_192_sva_dfm_1_1_enexo;
  assign act_port_reg_data_and_34_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_175_160_sva_dfm_1_1_enexo;
  assign act_port_reg_data_and_35_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_111_96_sva_dfm_1_1_enexo;
  assign act_port_reg_data_and_36_enex5 = act_port_reg_data_and_cse & reg_act_port_reg_data_143_128_sva_dfm_1_1_enexo;
  assign PECore_PushOutput_if_and_cse = PECoreRun_wen & and_dcpl_22;
  assign PECore_RunMac_if_and_cse = PECoreRun_wen & and_dcpl_25;
  assign while_if_and_6_cse = PECoreRun_wen & while_stage_0_10;
  assign PECore_RunMac_if_and_1_cse = PECoreRun_wen & (and_dcpl_28 | and_dcpl_305);
  assign while_if_and_7_cse = PECoreRun_wen & while_stage_0_9;
  assign PECore_RunMac_if_and_2_cse = PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & rva_in_reg_rw_sva_st_1_6)) & while_stage_0_8;
  assign while_if_and_8_cse = PECoreRun_wen & while_stage_0_8;
  assign weight_port_read_out_data_and_enex5 = PECoreRun_wen & (~((~ while_stage_0_8)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~ weight_mem_run_3_for_land_3_lpi_1_dfm_3))) & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_000000;
  assign weight_mem_run_3_for_aelse_and_cse = PECoreRun_wen & while_stage_0_7;
  assign and_536_itm = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  assign nor_413_itm = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | weight_mem_run_3_for_land_3_lpi_1_dfm_2);
  assign PECore_RunMac_if_and_3_cse = PECoreRun_wen & (~(rva_in_reg_rw_sva_st_1_5
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5))
      & while_stage_0_7;
  assign weight_mem_banks_read_1_read_data_and_8_cse = PECoreRun_wen & and_dcpl_44;
  assign input_mem_banks_read_1_read_data_and_2_enex5 = PECoreRun_wen & and_dcpl_44
      & reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  assign weight_mem_run_3_for_aelse_and_1_cse = PECoreRun_wen & while_stage_0_6;
  assign or_25_nl = and_679_cse | and_887_cse | and_889_cse | and_888_cse | and_890_cse
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]))
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | not_tmp_33;
  assign or_19_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7])) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | not_tmp_33;
  assign mux_10_nl = MUX_s_1_2_2(or_25_nl, or_19_nl, weight_mem_read_arbxbar_arbiters_next_7_6_sva);
  assign or_17_nl = (~ weight_mem_read_arbxbar_arbiters_next_7_6_sva) | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7])) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | not_tmp_33;
  assign mux_11_nl = MUX_s_1_2_2(mux_10_nl, or_17_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign or_15_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | nand_39_cse;
  assign mux_12_nl = MUX_s_1_2_2(mux_11_nl, or_15_nl, while_stage_0_5);
  assign or_13_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_run_3_for_land_7_lpi_1_dfm_1);
  assign mux_13_nl = MUX_s_1_2_2(mux_12_nl, or_13_nl, while_stage_0_6);
  assign weight_port_read_out_data_and_71_cse = PECoreRun_wen & weight_mem_run_3_for_land_7_lpi_1_dfm_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7 & fsm_output & mux_13_nl;
  assign weight_port_read_out_data_and_10_cse = PECoreRun_wen & (~(or_dcpl_218 |
      (~ weight_mem_run_3_for_land_2_lpi_1_dfm_2)));
  assign weight_port_read_out_data_and_18_cse = PECoreRun_wen & (~(or_dcpl_218 |
      (~ weight_mem_run_3_for_land_3_lpi_1_dfm_2)));
  assign weight_port_read_out_data_and_24_cse = PECoreRun_wen & (~((~ weight_mem_run_3_for_land_5_lpi_1_dfm_2)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7)));
  assign weight_port_read_out_data_and_32_cse = PECoreRun_wen & (~((~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7)));
  assign and_1010_cse = (((weight_read_addrs_7_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[2])) | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign nor_690_cse = ~((weight_read_addrs_7_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_339_nl = MUX_s_1_2_2((weight_read_addrs_7_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_7_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_7_lpi_1_dfm_3_2_0[0]);
  assign mux_340_cse = MUX_s_1_2_2(mux_339_nl, nor_690_cse, weight_read_addrs_7_lpi_1_dfm_3_2_0[2]);
  assign and_1018_cse = (mux_340_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign and_1019_cse = (and_1018_cse | or_dcpl_312 | weight_mem_run_3_for_5_and_156_itm_2
      | weight_mem_run_3_for_5_and_144_itm_1) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & PECoreRun_wen;
  assign and_1030_cse = (mux_340_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_port_read_out_data_5_7_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]), weight_port_read_out_data_5_7_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_316 , weight_mem_run_3_for_5_asn_318
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_320 , weight_mem_run_3_for_5_and_94_itm_1
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_and_96_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign nor_695_cse = ~((weight_read_addrs_5_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_349_nl = MUX_s_1_2_2((weight_read_addrs_5_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_5_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_5_lpi_1_dfm_3_2_0[0]);
  assign mux_350_nl = MUX_s_1_2_2(mux_349_nl, nor_695_cse, weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign and_1043_cse = (mux_350_nl | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign and_1044_cse = (and_1043_cse | weight_mem_run_3_for_5_and_96_itm_1 | weight_mem_run_3_for_5_and_95_itm_2
      | or_dcpl_345) & and_dcpl_719 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign weight_mem_run_3_for_5_and_81_nl = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_port_read_out_data_5_6_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]), weight_port_read_out_data_5_6_sva_dfm_1,
      {weight_mem_run_3_for_5_and_81_nl , weight_mem_run_3_for_5_asn_316 , weight_mem_run_3_for_5_asn_318
      , weight_mem_run_3_for_5_and_84_itm_1 , weight_mem_run_3_for_5_asn_320 , weight_mem_run_3_for_5_and_86_itm_2
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_asn_322 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign xor_7_cse = (weight_read_addrs_5_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_5_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign weight_port_read_out_data_5_5_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]), weight_port_read_out_data_5_5_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_316 , weight_mem_run_3_for_5_asn_318
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_320 , weight_mem_run_3_for_5_and_94_itm_1
      , weight_mem_run_3_for_5_and_79_itm_1 , weight_mem_run_3_for_5_and_96_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign and_1054_cse = (and_1043_cse | or_dcpl_355 | or_dcpl_345) & and_dcpl_719
      & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign weight_port_read_out_data_5_4_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]), weight_port_read_out_data_5_4_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_316 , weight_mem_run_3_for_5_asn_318
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_320 , weight_mem_run_3_for_5_and_86_itm_2
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_asn_322 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign and_1059_cse = (((xor_7_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2) | or_dcpl_350 | weight_mem_run_3_for_5_and_92_itm_2)
      & and_dcpl_719 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign weight_port_read_out_data_5_3_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]), weight_port_read_out_data_5_3_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_316 , weight_mem_run_3_for_5_asn_318
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_320 , weight_mem_run_3_for_5_and_94_itm_1
      , weight_mem_run_3_for_5_and_79_itm_1 , weight_mem_run_3_for_5_and_96_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_2_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]), weight_port_read_out_data_5_2_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_316 , weight_mem_run_3_for_5_asn_318
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_320 , weight_mem_run_3_for_5_and_86_itm_2
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_asn_322 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_1_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]), weight_port_read_out_data_5_1_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_316 , weight_mem_run_3_for_5_asn_318
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_320 , weight_mem_run_3_for_5_and_86_itm_2
      , weight_mem_run_3_for_5_and_79_itm_1 , weight_mem_run_3_for_5_and_96_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_0_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]),
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9, weight_port_read_out_data_5_0_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_316 , weight_mem_run_3_for_5_asn_318
      , weight_mem_run_3_for_5_and_92_itm_2 , weight_mem_run_3_for_5_asn_320 , weight_mem_run_3_for_5_and_94_itm_1
      , weight_mem_run_3_for_5_and_95_itm_2 , weight_mem_run_3_for_5_and_96_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_3_7_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]), weight_port_read_out_data_3_7_sva_dfm_1,
      {weight_mem_run_3_for_5_and_166 , weight_mem_run_3_for_5_asn_324 , weight_mem_run_3_for_5_asn_326
      , weight_mem_run_3_for_5_and_28_itm_1 , weight_mem_run_3_for_5_asn_328 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_31_itm_2 , weight_mem_run_3_for_5_asn_330 , (~
      weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign xor_13_cse = (weight_read_addrs_3_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_3_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_3_lpi_1_dfm_3_2_0[2]);
  assign and_1083_cse = (xor_13_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_port_read_out_data_3_6_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]), weight_port_read_out_data_3_6_sva_dfm_1,
      {weight_mem_run_3_for_5_and_166 , weight_mem_run_3_for_5_asn_324 , weight_mem_run_3_for_5_asn_326
      , weight_mem_run_3_for_5_and_20_itm_2 , weight_mem_run_3_for_5_asn_328 , weight_mem_run_3_for_5_and_22_itm_1
      , weight_mem_run_3_for_5_and_23_itm_1 , weight_mem_run_3_for_5_asn_330 , (~
      weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign weight_port_read_out_data_3_5_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]), weight_port_read_out_data_3_5_sva_dfm_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_73_cse , weight_mem_run_3_for_5_asn_324
      , weight_mem_run_3_for_5_asn_326 , weight_mem_run_3_for_5_and_20_itm_2 , weight_mem_run_3_for_5_asn_328
      , weight_mem_run_3_for_5_and_30_itm_2 , weight_mem_run_3_for_5_and_31_itm_2
      , weight_mem_run_3_for_5_asn_330 , (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign weight_mem_run_3_for_5_and_7_nl = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_port_read_out_data_3_4_sva_dfm_3 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]), weight_port_read_out_data_3_4_sva_dfm_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_73_cse , weight_mem_run_3_for_5_asn_324
      , weight_mem_run_3_for_5_asn_326 , weight_mem_run_3_for_5_and_20_itm_2 , weight_mem_run_3_for_5_asn_328
      , weight_mem_run_3_for_5_and_30_itm_2 , weight_mem_run_3_for_5_and_7_nl , weight_mem_run_3_for_5_and_8_itm_1
      , (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign weight_port_read_out_data_and_56_cse = PECoreRun_wen & (PECore_PushAxiRsp_and_2_cse
      | and_dcpl_375);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_101_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1 & while_stage_0_6 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_cse = PECoreRun_wen
      & or_tmp_60 & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_113_cse = PECoreRun_wen
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_2_lpi_1_dfm_1) & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_cse = PECoreRun_wen
      & and_dcpl_44 & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse = PECoreRun_wen & and_dcpl_44
      & weight_mem_run_3_for_land_1_lpi_1_dfm_2;
  assign and_706_cse = (Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign weight_read_addrs_and_7_enex5 = PECoreRun_wen & (and_dcpl_74 | (weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
      & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6])))) & and_882_cse &
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse = PECoreRun_wen & and_dcpl_81;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse
      & (reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo
      | reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1_enexo | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo);
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse = PECoreRun_wen & and_dcpl_83;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse
      & (reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1_enexo_1 | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2
      | reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1);
  assign while_if_and_11_cse = PECoreRun_wen & while_stage_0_5;
  assign weight_mem_read_arbxbar_arbiters_next_and_cse = PECoreRun_wen & fsm_output;
  assign weight_mem_read_arbxbar_arbiters_next_and_49_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((nor_226_cse & nor_227_cse & nor_228_cse & nor_229_cse) | or_dcpl_59);
  assign weight_mem_read_arbxbar_arbiters_next_and_55_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_107_cse | or_dcpl_59);
  assign weight_mem_read_arbxbar_arbiters_next_and_61_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_114_cse | or_dcpl_59);
  assign weight_mem_read_arbxbar_arbiters_next_and_67_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_121_cse | or_dcpl_59);
  assign weight_mem_read_arbxbar_arbiters_next_and_73_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_128_cse | or_dcpl_59);
  assign weight_mem_read_arbxbar_arbiters_next_and_79_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_135_cse | or_dcpl_59);
  assign weight_mem_read_arbxbar_arbiters_next_and_85_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_1_tmp) |
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4));
  assign weight_mem_read_arbxbar_arbiters_next_and_91_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & or_dcpl_68;
  assign weight_read_addrs_and_9_cse = PECoreRun_wen & (and_dcpl_147 | and_dcpl_146
      | and_dcpl_145 | and_dcpl_144 | and_dcpl_143 | and_dcpl_142 | and_dcpl_141
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | and_dcpl_140) & while_stage_0_4;
  assign weight_write_data_data_and_cse = PECoreRun_wen & and_dcpl_153 & ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7:6]!=2'b00));
  assign weight_write_data_data_and_24_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_25_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_26_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_27_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_28_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_29_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_30_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_31_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_addrs_and_enex5 = weight_write_data_data_and_cse & reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  assign weight_mem_write_arbxbar_xbar_for_1_for_and_cse = PECoreRun_wen & and_dcpl_153;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
      = PECoreRun_wen & and_dcpl_158;
  assign PECore_RunFSM_switch_lp_and_cse = PECoreRun_wen & while_stage_0_4;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 & and_dcpl_158;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 & and_dcpl_158;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12 & and_dcpl_158;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
      = PECoreRun_wen & (operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])) & and_dcpl_158;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_23_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_1_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign Arbiter_8U_Roundrobin_pick_1_and_15_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8
      & and_dcpl_158;
  assign Arbiter_8U_Roundrobin_pick_and_75_cse = PECoreRun_wen & (while_stage_0_4
      | and_dcpl_545) & fsm_output & or_dcpl_59;
  assign Arbiter_8U_Roundrobin_pick_1_and_22_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9
      & and_dcpl_158;
  assign Arbiter_8U_Roundrobin_pick_1_and_64_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15
      & and_dcpl_158;
  assign weight_write_data_data_and_8_cse = PECoreRun_wen & and_dcpl_194;
  assign weight_write_data_data_and_32_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_33_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_34_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_35_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_36_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_37_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_38_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_39_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  assign weight_write_addrs_and_2_enex5 = weight_write_data_data_and_8_cse & reg_pe_manager_base_input_enexo;
  assign rva_in_reg_rw_and_5_cse = PECoreRun_wen & while_stage_0_3;
  assign weight_read_addrs_and_28_enex5 = weight_write_data_data_and_8_cse & reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  assign state_and_cse = weight_mem_read_arbxbar_arbiters_next_and_cse & or_dcpl_135;
  assign and_1109_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & while_stage_0_3;
  assign pe_config_num_manager_and_cse = PECoreRun_wen & (~(or_dcpl_240 | or_dcpl_239
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~(PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])))));
  assign rva_in_reg_rw_and_6_cse = PECoreRun_wen & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign PECore_UpdateFSM_switch_lp_and_9_cse = PECoreRun_wen & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign or_220_cse = (state_2_1_sva!=2'b00) | state_0_sva;
  assign or_835_cse = (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_1884_cse = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  assign pe_config_UpdateManagerCounter_if_if_and_enex5 = PECoreRun_wen & reg_pe_config_num_output_enexo;
  assign PECore_DecodeAxiRead_switch_lp_and_cse = PECoreRun_wen & (~(or_dcpl_135
      | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
  assign PECore_DecodeAxiWrite_switch_lp_and_cse = PECoreRun_wen & (~ or_dcpl_239);
  assign or_228_cse_1 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
      | (~ while_stage_0_11);
  assign weight_mem_banks_load_store_for_else_and_cse = PECoreRun_wen & and_dcpl_43
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_101_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[55:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_101_nl);
  assign weight_mem_banks_load_store_for_else_and_6_cse = PECoreRun_wen & and_dcpl_43
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign or_713_tmp = ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]) & nor_260_cse)
      | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]) & and_dcpl_596) | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[2])
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]));
  assign weight_mem_banks_load_store_for_else_and_9_cse = PECoreRun_wen & while_stage_0_6
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign weight_mem_banks_load_store_for_else_and_10_cse = PECoreRun_wen & while_stage_0_6
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign or_231_cse = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]!=2'b00);
  assign weight_mem_banks_load_store_for_else_and_14_cse = PECoreRun_wen & and_dcpl_43
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1;
  assign weight_mem_banks_load_store_for_else_and_16_cse = PECoreRun_wen & and_dcpl_43
      & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]))
      & nor_260_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign weight_mem_banks_load_store_for_else_and_19_cse = PECoreRun_wen & and_dcpl_43
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[23:16]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl);
  assign weight_read_addrs_and_19_cse = PECoreRun_wen & and_dcpl_80;
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_103_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_99_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_75_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_24_cse
      = weight_mem_read_arbxbar_arbiters_next_and_cse & or_dcpl_59;
  assign weight_read_addrs_and_29_enex5 = weight_write_data_data_and_8_cse & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  assign operator_15_false_1_and_cse = PECoreRun_wen & (~(and_dcpl_544 | or_dcpl_59));
  assign PEManager_15U_PEManagerWrite_and_enex5 = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse & (~ PECore_DecodeAxiWrite_switch_lp_nor_tmp_1)
      & PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 & (~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1)) & while_stage_0_3 & reg_rva_in_reg_data_sva_1_enexo;
  assign pe_manager_num_input_and_cse = PECoreRun_wen & (~(or_dcpl_240 | or_dcpl_135
      | or_dcpl_275));
  assign pe_config_is_valid_and_cse = PECoreRun_wen & (~(PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1
      | PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (~ or_dcpl_135);
  assign nor_718_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:10]!=2'b00));
  assign and_1169_cse = (((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:2]==8'b00000000)
      & nor_718_cse & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:12]!=2'b00)))
      & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:14]!=2'b00))) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | (~(reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3))) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01)
      & rva_in_PopNB_mioi_return_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]==2'b00)
      & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & rva_in_reg_rw_and_6_cse;
  assign while_if_and_15_cse = PECoreRun_wen & and_dcpl_240;
  assign rva_in_reg_rw_and_7_cse = PECoreRun_wen & and_882_cse;
  assign while_if_and_16_cse = PECoreRun_wen & and_dcpl_245;
  assign or_261_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_122_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_74_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_79_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_1_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign weight_port_read_out_data_and_79_cse = PECoreRun_wen & and_dcpl_244 & (~
      rva_in_reg_rw_sva_st_1_8) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  assign input_mem_banks_read_read_data_and_9_cse = PECoreRun_wen & and_dcpl_267
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6) & input_read_req_valid_lpi_1_dfm_1_8;
  assign weight_port_read_out_data_and_95_enex5 = weight_port_read_out_data_and_79_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo;
  assign input_mem_banks_read_read_data_and_35_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  assign weight_port_read_out_data_and_96_enex5 = weight_port_read_out_data_and_79_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo;
  assign input_mem_banks_read_read_data_and_36_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo;
  assign weight_port_read_out_data_and_97_enex5 = weight_port_read_out_data_and_79_cse
      & reg_weight_port_read_out_data_0_2_sva_dfm_3_2_enexo;
  assign input_mem_banks_read_read_data_and_37_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_38_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse = PECoreRun_wen & and_dcpl_244
      & (~(rva_in_reg_rw_sva_st_1_8 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6))
      & (~(rva_in_reg_rw_sva_8 | input_read_req_valid_lpi_1_dfm_1_8)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  assign and_1197_cse = (PECore_UpdateFSM_switch_lp_equal_tmp_2_9 | (~ while_stage_0_11)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
      | (PECore_RunScale_PECore_RunScale_if_and_1_svs_8 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_8)))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & PECoreRun_wen & while_stage_0_10 & (PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8
      | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8));
  assign input_mem_banks_read_1_read_data_and_3_enex5 = PECoreRun_wen & ((PECore_RunMac_PECore_RunMac_if_and_svs_st_3
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5) | (and_dcpl_393 & input_read_req_valid_lpi_1_dfm_1_3 & and_882_cse))
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  assign or_286_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
      | and_713_cse;
  assign or_296_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp
      | and_715_cse;
  assign input_read_req_valid_and_1_cse = PECoreRun_wen & and_dcpl_267;
  assign PECore_DecodeAxiRead_switch_lp_and_7_cse = PECoreRun_wen & and_dcpl_284;
  assign rva_out_reg_data_and_24_cse = PECoreRun_wen & and_dcpl_284 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_8) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8)
      & (~(rva_in_reg_rw_sva_st_1_8 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8));
  assign rva_out_reg_data_and_93_enex5 = rva_out_reg_data_and_24_cse & reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_94_enex5 = rva_out_reg_data_and_24_cse & reg_rva_out_reg_data_23_17_sva_dfm_6_1_enexo;
  assign rva_out_reg_data_and_95_enex5 = rva_out_reg_data_and_24_cse & reg_rva_out_reg_data_15_9_sva_dfm_8_1_enexo;
  assign weight_port_read_out_data_and_98_enex5 = weight_port_read_out_data_and_79_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_3_2_enexo;
  assign rva_out_reg_data_and_96_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_97_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_98_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_99_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_100_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_3_1_enexo;
  assign weight_mem_run_3_for_weight_mem_run_3_for_and_4_cse = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & or_261_cse;
  assign and_1231_cse = (~((~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
      | (~ while_stage_0_10))) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9))
      & while_stage_0_11 & fsm_output & PECoreRun_wen;
  assign ProductSum_for_and_cse = PECoreRun_wen & and_dcpl_25 & (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
  assign weight_port_read_out_data_and_86_cse = PECoreRun_wen & and_dcpl_27 & (~
      rva_in_reg_rw_sva_st_1_7) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  assign and_1258_cse = (PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | PECore_UpdateFSM_switch_lp_equal_tmp_2_8)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & while_if_and_6_cse;
  assign PECore_RunScale_if_and_1_cse = PECoreRun_wen & and_dcpl_28;
  assign weight_mem_write_arbxbar_xbar_for_empty_and_enex5 = rva_in_reg_rw_and_7_cse
      & reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  assign and_301_cse = PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]);
  assign input_mem_banks_read_read_data_and_18_cse = PECoreRun_wen & and_dcpl_305
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5) & input_read_req_valid_lpi_1_dfm_1_7;
  assign input_mem_banks_read_read_data_and_39_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo;
  assign input_mem_banks_read_read_data_and_40_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_1;
  assign input_mem_banks_read_read_data_and_41_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_2;
  assign input_mem_banks_read_read_data_and_42_enex5 = input_mem_banks_read_read_data_and_18_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse = PECoreRun_wen & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6
      & while_stage_0_9 & and_dcpl_309 & and_dcpl_308;
  assign and_712_nl = input_read_req_valid_lpi_1_dfm_1_2 & not_tmp_182;
  assign mux_79_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2, and_712_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign input_mem_banks_read_1_read_data_and_4_enex5 = PECoreRun_wen & mux_79_nl
      & while_stage_0_4 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  assign input_read_req_valid_and_2_cse = PECoreRun_wen & and_dcpl_305;
  assign PECore_DecodeAxiRead_switch_lp_and_11_cse = PECoreRun_wen & and_dcpl_305
      & and_dcpl_308;
  assign rva_out_reg_data_and_34_cse = PECoreRun_wen & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 | rva_in_reg_rw_sva_st_1_7))
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_7) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6
      & while_stage_0_9 & and_dcpl_309 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5)
      & (~(rva_in_reg_rw_sva_7 | input_read_req_valid_lpi_1_dfm_1_7));
  assign rva_out_reg_data_and_101_enex5 = rva_out_reg_data_and_34_cse & reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_102_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_103_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo;
  assign input_mem_banks_read_read_data_and_27_enex5 = PECoreRun_wen & and_dcpl_325
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4) & input_read_req_valid_lpi_1_dfm_1_6
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0_enexo;
  assign PECore_RunMac_if_and_6_cse = PECoreRun_wen & and_604_cse;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse = PECoreRun_wen & and_dcpl_30
      & (~(rva_in_reg_rw_sva_st_1_6 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4))
      & (~(rva_in_reg_rw_sva_6 | input_read_req_valid_lpi_1_dfm_1_6)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
  assign nor_308_nl = ~((~ input_read_req_valid_lpi_1_dfm_1_1) | reg_rva_in_reg_rw_sva_st_1_1_cse);
  assign mux_80_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_3_1, nor_308_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign input_mem_banks_read_1_read_data_and_5_enex5 = PECoreRun_wen & mux_80_nl
      & while_stage_0_3 & (reg_input_mem_banks_bank_a_23_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_131_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_15_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_76_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_126_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_73_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_252_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_96_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_77_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_127_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_22_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_140_sva_dfm_2_enexo
      | reg_input_read_addrs_sva_1_1_enexo | reg_input_mem_banks_bank_a_157_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_183_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_11_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_236_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_64_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_109_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_195_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_17_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_228_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_147_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_32_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_184_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_9_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_162_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_188_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_14_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_35_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_207_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_49_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_238_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_130_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_53_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_179_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_106_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_70_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_185_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_113_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_90_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_197_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_146_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_88_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_85_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_108_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_112_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_7_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_255_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_221_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_227_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_33_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_192_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_142_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_141_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_151_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_41_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_61_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_167_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_119_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_115_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_63_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_71_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_229_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_103_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_143_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_59_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_189_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_204_sva_dfm_2_enexo | reg_input_mem_banks_read_read_data_sva_1_enexo
      | reg_input_mem_banks_bank_a_166_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_31_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_214_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_220_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_27_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_163_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_139_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_78_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_249_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_99_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_8_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_26_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_100_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_20_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_226_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_79_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_134_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_161_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_82_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_24_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_36_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_75_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_6_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_232_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_187_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_218_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_239_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_42_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_124_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_152_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_164_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_180_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_3_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_107_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_39_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_186_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_45_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_125_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_198_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_87_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_196_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_160_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_171_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_135_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_149_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_60_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_80_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_170_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_159_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_81_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_104_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_84_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_194_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_136_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_118_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_40_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_243_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_148_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_177_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_91_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_16_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_66_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_237_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_138_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_219_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_213_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_199_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_230_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_117_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_47_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_244_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_231_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_172_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_240_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_34_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_191_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_173_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_121_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_245_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_105_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_181_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_69_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_89_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_169_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_193_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_5_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_200_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_212_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_137_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_21_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_58_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_12_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_1_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_174_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_155_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_211_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_18_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_190_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_116_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_97_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_54_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_29_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_122_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_55_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_224_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_206_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_13_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_253_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_201_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_94_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_37_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_28_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_132_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_92_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_215_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_62_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_38_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_223_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_242_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_233_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_154_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_235_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_72_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_250_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_129_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_234_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_98_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_10_sva_dfm_2_enexo
      | reg_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1_enexo
      | reg_input_mem_banks_bank_a_44_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_30_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_133_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_225_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_68_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_210_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_251_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_202_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_247_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_182_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_175_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_145_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_123_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_86_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_52_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_48_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_83_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_95_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_102_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_222_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_114_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_246_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_110_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_153_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_2_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_65_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_128_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_209_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_0_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_25_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_46_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_217_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_205_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_248_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_57_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_216_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_74_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_120_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_93_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_168_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_4_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_50_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_254_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_101_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_165_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_176_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_203_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_43_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_208_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_144_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_156_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_67_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_178_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_56_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_111_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_158_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_150_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_19_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_241_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_51_sva_dfm_2_enexo);
  assign input_read_req_valid_and_3_cse = PECoreRun_wen & and_dcpl_325;
  assign PECore_DecodeAxiRead_switch_lp_and_15_cse = PECoreRun_wen & and_dcpl_337;
  assign rva_out_reg_data_and_42_cse = PECoreRun_wen & and_dcpl_337 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5
      & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6)
      & (~(rva_in_reg_rw_sva_st_1_6 | PECore_DecodeAxiRead_switch_lp_nor_tmp_6));
  assign rva_out_reg_data_and_104_enex5 = rva_out_reg_data_and_42_cse & reg_rva_out_reg_data_30_25_sva_dfm_4_enexo;
  assign rva_out_reg_data_and_105_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_106_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo;
  assign PECore_RunScale_if_and_2_cse = PECoreRun_wen & while_stage_0_8 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6);
  assign or_898_cse = (state_2_1_sva[1]) | state_0_sva;
  assign nor_744_nl = ~((state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt));
  assign mux_365_cse = MUX_s_1_2_2(nor_744_nl, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_898_cse);
  assign nand_247_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b11));
  assign nand_248_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2:0]==3'b111));
  assign nor_776_nl = ~((state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign nor_777_nl = ~((~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign mux_387_cse = MUX_s_1_2_2(nor_776_nl, nor_777_nl, or_898_cse);
  assign or_977_nl = (state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[0]));
  assign or_975_nl = (~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[0]));
  assign mux_389_cse = MUX_s_1_2_2(or_977_nl, or_975_nl, or_898_cse);
  assign nand_250_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3:0]==4'b1111));
  assign or_1015_nl = (state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[2]));
  assign or_1013_nl = (~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[2]));
  assign mux_403_cse = MUX_s_1_2_2(or_1015_nl, or_1013_nl, or_898_cse);
  assign or_1054_nl = (state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[1]));
  assign or_1052_nl = (~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[1]));
  assign mux_415_cse = MUX_s_1_2_2(or_1054_nl, or_1052_nl, or_898_cse);
  assign nor_816_nl = ~((state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[1])));
  assign nor_817_nl = ~((~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[1])));
  assign mux_417_cse = MUX_s_1_2_2(nor_816_nl, nor_817_nl, or_898_cse);
  assign nand_254_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4:0]==5'b11111));
  assign nand_262_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5:0]==6'b111111));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse = PECoreRun_wen & and_dcpl_350
      & and_dcpl_349 & while_stage_0_7 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign input_mem_banks_read_read_data_and_28_enex5 = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      & (~ rva_in_reg_rw_sva_st_1_5) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  assign input_read_req_valid_and_4_cse = PECoreRun_wen & and_dcpl_357;
  assign PECore_DecodeAxiRead_switch_lp_and_19_cse = PECoreRun_wen & and_dcpl_350
      & (~ rva_in_reg_rw_sva_st_1_5) & PECore_PushAxiRsp_and_2_cse & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign rva_out_reg_data_and_50_enex5 = PECoreRun_wen & and_dcpl_350 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5)
      & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5))
      & (~ rva_in_reg_rw_sva_st_1_5) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      & reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_1_enexo;
  assign rva_out_reg_data_and_51_cse = PECoreRun_wen & (~(rva_in_reg_rw_sva_5 & rva_in_reg_rw_sva_st_1_5))
      & PECore_PushAxiRsp_and_2_cse;
  assign and_1792_cse = (~(((~(rva_in_reg_rw_sva_6 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      | (~ while_stage_0_8) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)) | rva_in_reg_rw_sva_st_1_5)
      & rva_in_reg_rw_sva_5)) & PECore_PushAxiRsp_and_2_cse & PECoreRun_wen;
  assign PECore_RunScale_if_and_3_cse = PECoreRun_wen & and_dcpl_375;
  assign or_317_nl = (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      | (~ reg_rva_in_PopNB_mioi_iswt0_cse);
  assign or_315_nl = reg_rva_in_reg_rw_sva_st_1_1_cse | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_86_nl = MUX_s_1_2_2(or_317_nl, or_315_nl, while_stage_0_3);
  assign or_314_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      | reg_rva_in_reg_rw_sva_2_cse;
  assign mux_87_nl = MUX_s_1_2_2(mux_86_nl, or_314_nl, while_stage_0_4);
  assign or_313_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      | rva_in_reg_rw_sva_3;
  assign mux_88_nl = MUX_s_1_2_2(mux_87_nl, or_313_nl, while_stage_0_5);
  assign or_312_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | rva_in_reg_rw_sva_4;
  assign mux_89_nl = MUX_s_1_2_2(mux_88_nl, or_312_nl, while_stage_0_6);
  assign or_305_nl = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      | rva_in_reg_rw_sva_5;
  assign mux_85_cse = MUX_s_1_2_2(mux_89_nl, or_305_nl, while_stage_0_7);
  assign rva_out_reg_data_and_56_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & mux_85_cse;
  assign and_1801_cse = mux_85_cse & and_dcpl_30 & (~ rva_in_reg_rw_sva_6) & weight_mem_read_arbxbar_arbiters_next_and_cse;
  assign PECore_PushAxiRsp_and_2_cse = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7;
  assign mux_70_nl = MUX_s_1_2_2((~ or_tmp_84), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign rva_out_reg_data_and_61_cse = PECoreRun_wen & mux_70_nl & and_dcpl_43;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse = PECoreRun_wen & (~ rva_in_reg_rw_sva_4)
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 & and_dcpl_43 & (~(rva_in_reg_rw_sva_st_1_4
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2));
  assign mux_91_nl = MUX_s_1_2_2((~ weight_mem_run_3_for_land_4_lpi_1_dfm_1), rva_in_reg_rw_sva_4,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_92_nl = MUX_s_1_2_2(mux_91_nl, or_38_cse, or_tmp_2);
  assign PECore_DecodeAxiRead_switch_lp_and_23_cse = PECoreRun_wen & (~ mux_92_nl)
      & while_stage_0_6;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_23_cse = PECoreRun_wen & and_dcpl_393
      & (~(input_read_req_valid_lpi_1_dfm_1_3 | rva_in_reg_rw_sva_3)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_713_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5;
  assign nand_39_cse = ~(or_286_cse & PECore_RunFSM_switch_lp_equal_tmp_1_2);
  assign and_715_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1;
  assign nor_284_nl = ~(rva_in_reg_rw_sva_3 | input_read_req_valid_lpi_1_dfm_1_3
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 | rva_in_reg_rw_sva_st_1_3);
  assign mux_96_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, nor_284_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign PECore_DecodeAxiRead_switch_lp_and_27_cse = PECoreRun_wen & mux_96_nl &
      while_stage_0_5;
  assign rva_out_reg_data_and_62_cse = PECoreRun_wen & and_dcpl_406 & (~(rva_in_reg_rw_sva_3
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_3)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3
      | rva_in_reg_rw_sva_st_1_3)) & and_882_cse;
  assign rva_out_reg_data_and_107_enex5 = rva_out_reg_data_and_62_cse & reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_108_enex5 = rva_out_reg_data_and_62_cse & reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_109_enex5 = rva_out_reg_data_and_62_cse & reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_65_cse = PECoreRun_wen & and_dcpl_406 & (~ rva_in_reg_rw_sva_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign rva_out_reg_data_and_110_enex5 = rva_out_reg_data_and_65_cse & reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_111_enex5 = rva_out_reg_data_and_65_cse & reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_112_enex5 = rva_out_reg_data_and_65_cse & reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_113_enex5 = rva_out_reg_data_and_65_cse & reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_114_enex5 = rva_out_reg_data_and_65_cse & reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_28_cse = PECoreRun_wen & and_dcpl_417
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 & and_dcpl_153;
  assign PECore_DecodeAxiRead_switch_lp_and_31_cse = PECoreRun_wen & and_dcpl_417
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign rva_out_reg_data_and_70_cse = PECoreRun_wen & not_tmp_182 & (~(input_read_req_valid_lpi_1_dfm_1_2
      | reg_rva_in_reg_rw_sva_2_cse | PECore_DecodeAxiRead_switch_lp_nor_tmp_2))
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2)
      & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2) & and_dcpl_153;
  assign rva_out_reg_data_and_115_enex5 = rva_out_reg_data_and_70_cse & reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  assign rva_out_reg_data_and_116_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_117_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_118_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_119_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_120_enex5 = PECore_DecodeAxiRead_switch_lp_and_31_cse
      & reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_33_cse = PECoreRun_wen & mux_tmp_97
      & and_dcpl_435;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse = PECoreRun_wen & (~ reg_rva_in_reg_rw_sva_st_1_1_cse)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_switch_lp_and_35_cse = PECoreRun_wen & and_dcpl_435;
  assign rva_out_reg_data_and_78_enex5 = PECoreRun_wen & (~(input_read_req_valid_lpi_1_dfm_1_1
      | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[0])))
      & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[3:1]==3'b010)
      & and_dcpl_441 & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_121_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_122_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_123_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_124_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_125_enex5 = PECore_DecodeAxiRead_switch_lp_and_35_cse
      & reg_rva_out_reg_data_55_48_sva_dfm_1_1_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse = PECoreRun_wen & mux_tmp_97
      & and_dcpl_434 & (~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1) &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse = PECoreRun_wen & and_dcpl_207
      & and_dcpl_209 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse = PECoreRun_wen & and_dcpl_297
      & (~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])))
      & nand_31_cse;
  assign rva_out_reg_data_and_85_cse = PECoreRun_wen & (or_dcpl_141 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]!=2'b10))
      & and_dcpl_245;
  assign or_708_cse = ((Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 |
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse) & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1)
      | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp;
  assign and_882_cse = while_stage_0_5 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign and_522_cse = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
      & while_stage_0_12 & (~ rva_in_reg_rw_sva_st_1_10);
  assign weight_mem_run_3_for_5_and_177_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_175_cse = reg_weight_mem_run_3_for_5_and_162_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_176_cse = reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_178_cse = reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_182_cse = reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_189_cse = reg_weight_mem_run_3_for_5_and_168_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_197_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_196_cse = reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_203_cse = reg_weight_mem_run_3_for_5_and_166_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_port_read_out_data_7_6_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]), weight_port_read_out_data_7_6_sva_dfm_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_308 , weight_mem_run_3_for_5_asn_310
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_312 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_159_itm_1 , weight_mem_run_3_for_5_asn_314 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_7_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]), weight_port_read_out_data_7_7_sva_dfm_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_308 , weight_mem_run_3_for_5_asn_310
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_312 , weight_mem_run_3_for_5_and_158_itm_1
      , weight_mem_run_3_for_5_and_159_itm_1 , weight_mem_run_3_for_5_asn_314 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_4_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]), weight_port_read_out_data_7_4_sva_dfm_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_308 , weight_mem_run_3_for_5_asn_310
      , weight_mem_run_3_for_5_and_132_itm_1 , weight_mem_run_3_for_5_asn_312 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_159_itm_1 , weight_mem_run_3_for_5_asn_314 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_5_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]), weight_port_read_out_data_7_5_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_308 , weight_mem_run_3_for_5_asn_310
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_312 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_159_itm_1 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_2_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]), weight_port_read_out_data_7_2_sva_dfm_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_308 , weight_mem_run_3_for_5_asn_310
      , weight_mem_run_3_for_5_and_132_itm_1 , weight_mem_run_3_for_5_asn_312 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_159_itm_1 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_3_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]), weight_port_read_out_data_7_3_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_308 , weight_mem_run_3_for_5_asn_310
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_312 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_159_itm_1 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_0_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]),
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9, weight_port_read_out_data_7_0_sva_dfm_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_308 , weight_mem_run_3_for_5_asn_310
      , weight_mem_run_3_for_5_and_132_itm_1 , weight_mem_run_3_for_5_asn_312 , weight_mem_run_3_for_5_and_150_itm_2
      , weight_mem_run_3_for_5_and_103_itm_2 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_1_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]), weight_port_read_out_data_7_1_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_308 , weight_mem_run_3_for_5_asn_310
      , weight_mem_run_3_for_5_and_132_itm_1 , weight_mem_run_3_for_5_asn_312 , weight_mem_run_3_for_5_and_158_itm_1
      , weight_mem_run_3_for_5_and_159_itm_1 , weight_mem_run_3_for_5_and_144_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      | (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1:0]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]) & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_927_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_dcpl_302);
  assign and_928_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56 & (~ or_dcpl_302);
  assign and_929_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse & (~ or_dcpl_302);
  assign and_930_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      & (~ or_dcpl_302);
  assign and_931_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1
      & (~ or_dcpl_302);
  assign and_932_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1
      & (~ or_dcpl_302);
  assign and_933_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1
      & (~ or_dcpl_302);
  assign nor_426_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl_302);
  assign and_937_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56 & (~ or_dcpl_303);
  assign and_938_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse & (~ or_dcpl_303);
  assign and_939_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      & (~ or_dcpl_303);
  assign and_940_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1
      & (~ or_dcpl_303);
  assign and_941_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1
      & (~ or_dcpl_303);
  assign and_942_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1
      & (~ or_dcpl_303);
  assign nor_427_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl_303);
  assign PECore_PushAxiRsp_if_else_mux_13_mx0w2 = MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1);
  assign while_and_24_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign while_and_23_cse = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1_1
      = ~((weight_read_addrs_3_lpi_1_dfm_2_2_0!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign Arbiter_8U_Roundrobin_pick_nand_56_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1)
      & and_dcpl_80)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_36_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1
      & and_dcpl_80;
  assign weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_56_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_56_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_56_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_56_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_56_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0 = weight_mem_read_arbxbar_arbiters_next_7_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_7_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_56_cse , Arbiter_8U_Roundrobin_pick_and_36_cse});
  assign weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_80);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign Arbiter_8U_Roundrobin_pick_nand_44_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)
      & and_dcpl_80)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_30_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1
      & and_dcpl_80;
  assign weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_44_cse , Arbiter_8U_Roundrobin_pick_and_30_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_44_cse , Arbiter_8U_Roundrobin_pick_and_30_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_44_cse , Arbiter_8U_Roundrobin_pick_and_30_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_44_cse , Arbiter_8U_Roundrobin_pick_and_30_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_44_cse , Arbiter_8U_Roundrobin_pick_and_30_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0 = weight_mem_read_arbxbar_arbiters_next_6_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_6_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_44_cse , Arbiter_8U_Roundrobin_pick_and_30_cse});
  assign weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_80);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign Arbiter_8U_Roundrobin_pick_nand_32_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1)
      & and_dcpl_80)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_24_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1
      & and_dcpl_80;
  assign weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_32_cse , Arbiter_8U_Roundrobin_pick_and_24_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_32_cse , Arbiter_8U_Roundrobin_pick_and_24_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_39_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_39_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_32_cse , Arbiter_8U_Roundrobin_pick_and_24_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_38_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_38_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_32_cse , Arbiter_8U_Roundrobin_pick_and_24_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_37_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_37_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_32_cse , Arbiter_8U_Roundrobin_pick_and_24_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_32_cse , Arbiter_8U_Roundrobin_pick_and_24_cse});
  assign weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_80);
  assign Arbiter_8U_Roundrobin_pick_nand_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1)
      & and_dcpl_80)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_38_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1
      & and_dcpl_80;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_74_nl = weight_mem_read_arbxbar_arbiters_next_4_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_74_nl,
      weight_mem_read_arbxbar_arbiters_next_4_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_nl = weight_mem_read_arbxbar_arbiters_next_4_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_75_nl,
      weight_mem_read_arbxbar_arbiters_next_4_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_76_nl = weight_mem_read_arbxbar_arbiters_next_4_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_76_nl,
      weight_mem_read_arbxbar_arbiters_next_4_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_77_nl = weight_mem_read_arbxbar_arbiters_next_4_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_77_nl,
      weight_mem_read_arbxbar_arbiters_next_4_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_nl = weight_mem_read_arbxbar_arbiters_next_4_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_78_nl,
      weight_mem_read_arbxbar_arbiters_next_4_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_79_nl = weight_mem_read_arbxbar_arbiters_next_4_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_79_nl,
      weight_mem_read_arbxbar_arbiters_next_4_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_38_cse});
  assign weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_80);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign Arbiter_8U_Roundrobin_pick_nand_20_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1)
      & and_dcpl_80)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_18_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1
      & and_dcpl_80;
  assign weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_18_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_18_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_18_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_18_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_18_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_20_cse , Arbiter_8U_Roundrobin_pick_and_18_cse});
  assign weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_80);
  assign Arbiter_8U_Roundrobin_pick_nand_69_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1)
      & and_dcpl_80)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_50_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1
      & and_dcpl_80;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl = weight_mem_read_arbxbar_arbiters_next_2_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_86_nl,
      weight_mem_read_arbxbar_arbiters_next_2_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_50_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl = weight_mem_read_arbxbar_arbiters_next_2_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_87_nl,
      weight_mem_read_arbxbar_arbiters_next_2_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_50_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl = weight_mem_read_arbxbar_arbiters_next_2_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_88_nl,
      weight_mem_read_arbxbar_arbiters_next_2_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_50_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl = weight_mem_read_arbxbar_arbiters_next_2_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_89_nl,
      weight_mem_read_arbxbar_arbiters_next_2_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_50_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl = weight_mem_read_arbxbar_arbiters_next_2_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_90_nl,
      weight_mem_read_arbxbar_arbiters_next_2_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_50_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl = weight_mem_read_arbxbar_arbiters_next_2_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_91_nl,
      weight_mem_read_arbxbar_arbiters_next_2_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_50_cse});
  assign weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_80);
  assign Arbiter_8U_Roundrobin_pick_nand_81_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1)
      & and_dcpl_80)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_62_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1
      & and_dcpl_80;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_92_nl = weight_mem_read_arbxbar_arbiters_next_1_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_92_nl,
      weight_mem_read_arbxbar_arbiters_next_1_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_81_cse , Arbiter_8U_Roundrobin_pick_and_62_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl = weight_mem_read_arbxbar_arbiters_next_1_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_93_nl,
      weight_mem_read_arbxbar_arbiters_next_1_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_81_cse , Arbiter_8U_Roundrobin_pick_and_62_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl = weight_mem_read_arbxbar_arbiters_next_1_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_94_nl,
      weight_mem_read_arbxbar_arbiters_next_1_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_81_cse , Arbiter_8U_Roundrobin_pick_and_62_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_95_nl = weight_mem_read_arbxbar_arbiters_next_1_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_95_nl,
      weight_mem_read_arbxbar_arbiters_next_1_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_81_cse , Arbiter_8U_Roundrobin_pick_and_62_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl = weight_mem_read_arbxbar_arbiters_next_1_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_96_nl,
      weight_mem_read_arbxbar_arbiters_next_1_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_81_cse , Arbiter_8U_Roundrobin_pick_and_62_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_97_nl,
      weight_mem_read_arbxbar_arbiters_next_1_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_81_cse , Arbiter_8U_Roundrobin_pick_and_62_cse});
  assign weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_80);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign Arbiter_8U_Roundrobin_pick_nand_8_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1)
      & and_dcpl_80)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_12_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1
      & and_dcpl_80;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_12_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_4_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_4_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_12_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl = weight_mem_read_arbxbar_arbiters_next_0_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl,
      weight_mem_read_arbxbar_arbiters_next_0_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_12_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_2_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_2_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_12_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1,
      {and_882_cse , Arbiter_8U_Roundrobin_pick_nand_8_cse , Arbiter_8U_Roundrobin_pick_and_12_cse});
  assign weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_80);
  assign pe_manager_base_weight_sva_mx1_3_0 = MUX_v_4_2_2((pe_manager_base_weight_sva[3:0]),
      (pe_manager_base_weight_sva_dfm_3_1[3:0]), while_stage_0_5);
  assign pe_manager_base_weight_sva_mx2 = MUX_v_15_2_2(pe_manager_base_weight_sva,
      pe_manager_base_weight_sva_dfm_3_1, while_stage_0_5);
  assign nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000001;
  assign PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_1_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000001;
  assign operator_15_false_acc_nl = nl_operator_15_false_acc_nl[13:0];
  assign weight_read_addrs_2_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000011;
  assign PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_3_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_1_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:2])}) + 13'b0000000000001;
  assign operator_15_false_acc_1_nl = nl_operator_15_false_acc_1_nl[12:0];
  assign weight_read_addrs_4_14_2_lpi_1_dfm_1_1 = MUX_v_13_2_2(13'b0000000000000,
      operator_15_false_acc_1_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000101;
  assign PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_5_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_2_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000011;
  assign operator_15_false_acc_2_nl = nl_operator_15_false_acc_2_nl[13:0];
  assign weight_read_addrs_6_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_2_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000111;
  assign PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_7_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112, and_dcpl_544);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97, and_107_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82, and_114_cse);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_23_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67, and_121_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52, and_128_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37, and_135_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign and_628_nl = (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1])))
      & (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])));
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22, and_628_nl);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl
      & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_1_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_1_tmp = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7, and_142_cse);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp = Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1 = (state_2_1_sva[0]) & (~((state_2_1_sva[1])
      | state_0_sva));
  assign state_mux_1_cse = MUX_v_2_2_2(state_2_1_sva, state_2_1_sva_dfm_1, while_stage_0_3);
  assign state_0_sva_mx1 = MUX_s_1_2_2(PECore_UpdateFSM_next_state_0_lpi_1_dfm_4,
      state_0_sva, or_dcpl_228);
  assign pe_config_manager_counter_sva_mx1 = MUX_v_4_2_2(pe_config_manager_counter_sva,
      pe_config_manager_counter_sva_dfm_3_1, and_1109_cse);
  assign PECore_PushOutput_PECore_PushOutput_if_and_svs_1 = (state_mux_1_cse[1])
      & (~((state_mux_1_cse[0]) | state_0_sva_mx1));
  assign PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1 = ~(PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_220_cse);
  assign pe_config_input_counter_and_cse = while_if_and_tmp_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign nl_operator_8_false_acc_nl = pe_config_input_counter_sva + 8'b00000001;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[7:0];
  assign pe_config_UpdateInputCounter_not_nl = ~ pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl = MUX_v_8_2_2(8'b00000000,
      operator_8_false_acc_nl, pe_config_UpdateInputCounter_not_nl);
  assign pe_config_input_counter_nand_nl = ~(while_stage_0_3 & (~((~(PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1129_cse_1)));
  assign while_and_4_nl = PECore_UpdateFSM_switch_lp_equal_tmp_3_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign pe_config_input_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_input_counter_sva,
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl, pe_config_input_counter_sva_dfm_1,
      {pe_config_input_counter_nand_nl , while_and_4_nl , pe_config_input_counter_and_cse});
  assign nl_operator_8_false_1_acc_nl = pe_config_output_counter_sva + 8'b00000001;
  assign operator_8_false_1_acc_nl = nl_operator_8_false_1_acc_nl[7:0];
  assign pe_config_UpdateManagerCounter_if_not_9_nl = ~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl
      = MUX_v_8_2_2(8'b00000000, operator_8_false_1_acc_nl, pe_config_UpdateManagerCounter_if_not_9_nl);
  assign pe_config_output_counter_nand_nl = ~(while_stage_0_3 & (~((~(and_1884_cse
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1129_cse_1)));
  assign while_and_63_nl = and_1884_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign pe_config_output_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_output_counter_sva,
      pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl,
      pe_config_output_counter_sva_dfm_1, {pe_config_output_counter_nand_nl , while_and_63_nl
      , pe_config_input_counter_and_cse});
  assign and_604_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_if_and_2_m1c = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & and_604_cse;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl
      = pe_config_is_zero_first_sva & (~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1);
  assign while_if_or_nl = (~((~((~ PECore_UpdateFSM_switch_lp_equal_tmp_5_1) & and_604_cse))
      & while_stage_0_3)) | ((~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1)
      & while_if_and_2_m1c);
  assign while_if_and_4_nl = pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
      & while_if_and_2_m1c;
  assign pe_config_is_zero_first_sva_mx1 = MUX1HOT_s_1_3_2(while_if_mux_19_itm_1,
      pe_config_is_zero_first_sva, pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl,
      {and_dcpl_194 , while_if_or_nl , while_if_and_4_nl});
  assign PECore_UpdateFSM_switch_lp_equal_tmp_6 = state_0_sva_mx1 & (state_mux_1_cse==2'b00);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1 = (state_mux_1_cse[0])
      & (~((state_mux_1_cse[1]) | state_0_sva_mx1));
  assign pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1
      = ~((pe_config_manager_counter_sva_mx1 != (operator_4_false_acc_sdt_sva_1[3:0]))
      | (operator_4_false_acc_sdt_sva_1[4]));
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0110);
  assign PECore_UpdateFSM_switch_lp_not_16_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_10;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_nl
      = MUX_v_16_2_2(16'b0000000000000000, act_port_reg_data_79_64_sva_dfm_1_1, PECore_UpdateFSM_switch_lp_not_16_nl);
  assign or_452_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
      | (~ while_stage_0_12);
  assign act_port_reg_data_79_64_sva_mx1 = MUX_v_16_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_nl,
      act_port_reg_data_79_64_sva, or_452_nl);
  assign weight_mem_run_3_for_land_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_103_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1);
  assign weight_mem_run_3_for_land_6_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_75_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_99_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_111_tmp | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1);
  assign weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp);
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  assign weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6,
      or_dcpl_227);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0,
      or_dcpl_227);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5,
      or_dcpl_227);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1,
      or_dcpl_227);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4,
      or_dcpl_227);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2,
      or_dcpl_227);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3,
      or_dcpl_227);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0101);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b111)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b110)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b100)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b010)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b001)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_111_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
  assign PECore_UpdateFSM_switch_lp_not_26_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_nl
      = MUX_v_16_2_2(16'b0000000000000000, act_port_reg_data_15_0_sva_dfm_1_1, PECore_UpdateFSM_switch_lp_not_26_nl);
  assign act_port_reg_data_15_0_sva_mx1 = MUX_v_16_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_nl,
      act_port_reg_data_15_0_sva, or_228_cse_1);
  assign PECore_UpdateFSM_switch_lp_not_27_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_nl
      = MUX_v_16_2_2(16'b0000000000000000, act_port_reg_data_47_32_sva_dfm_1_1, PECore_UpdateFSM_switch_lp_not_27_nl);
  assign act_port_reg_data_47_32_sva_mx1 = MUX_v_16_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_nl,
      act_port_reg_data_47_32_sva, or_228_cse_1);
  assign PECore_UpdateFSM_switch_lp_not_28_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_nl
      = MUX_v_16_2_2(16'b0000000000000000, act_port_reg_data_111_96_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_28_nl);
  assign act_port_reg_data_111_96_sva_mx1 = MUX_v_16_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_nl,
      act_port_reg_data_111_96_sva, or_228_cse_1);
  assign PECore_UpdateFSM_switch_lp_not_29_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_11_nl
      = MUX_v_16_2_2(16'b0000000000000000, act_port_reg_data_143_128_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_29_nl);
  assign act_port_reg_data_143_128_sva_mx1 = MUX_v_16_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_11_nl,
      act_port_reg_data_143_128_sva, or_228_cse_1);
  assign PECore_UpdateFSM_switch_lp_not_30_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_10_nl
      = MUX_v_16_2_2(16'b0000000000000000, act_port_reg_data_175_160_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_30_nl);
  assign act_port_reg_data_175_160_sva_mx1 = MUX_v_16_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_10_nl,
      act_port_reg_data_175_160_sva, or_228_cse_1);
  assign PECore_UpdateFSM_switch_lp_not_31_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_9_nl
      = MUX_v_16_2_2(16'b0000000000000000, act_port_reg_data_207_192_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_31_nl);
  assign act_port_reg_data_207_192_sva_mx1 = MUX_v_16_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_9_nl,
      act_port_reg_data_207_192_sva, or_228_cse_1);
  assign PECore_UpdateFSM_switch_lp_not_25_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl
      = MUX_v_16_2_2(16'b0000000000000000, act_port_reg_data_239_224_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_25_nl);
  assign act_port_reg_data_239_224_sva_mx1 = MUX_v_16_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl,
      act_port_reg_data_239_224_sva, or_228_cse_1);
  assign weight_mem_run_3_for_land_1_lpi_1_dfm_1_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_23_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1 = MUX_v_3_2_2(3'b000,
      (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0]), weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_1_tmp = MUX_s_1_8_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_1_tmp
      | (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp));
  assign while_or_2_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_2_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_100_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_2_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_101_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_tmp_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_0_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_0_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_2_nl
      , while_and_100_nl , while_and_101_nl});
  assign while_or_3_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_3_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_1_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_104_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_3_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_105_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_1_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_1_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_1_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_3_nl
      , while_and_104_nl , while_and_105_nl});
  assign while_or_4_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_4_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_2_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_108_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_4_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_109_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_2_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_2_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_2_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_4_nl
      , while_and_108_nl , while_and_109_nl});
  assign while_or_5_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_5_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_3_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_112_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_5_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_113_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_3_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_3_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_3_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_5_nl
      , while_and_112_nl , while_and_113_nl});
  assign while_or_6_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_6_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_4_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_116_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_6_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_117_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_4_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_4_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_4_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_6_nl
      , while_and_116_nl , while_and_117_nl});
  assign while_or_7_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_7_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_5_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_120_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_7_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_121_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_5_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_5_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_5_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_7_nl
      , while_and_120_nl , while_and_121_nl});
  assign while_or_8_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_8_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_6_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_124_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_8_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_125_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_6_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_6_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_6_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_8_nl
      , while_and_124_nl , while_and_125_nl});
  assign while_or_9_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_9_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_7_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_128_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_9_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_129_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_7_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_7_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_7_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_9_nl
      , while_and_128_nl , while_and_129_nl});
  assign while_or_10_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_10_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_8_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_132_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_10_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_133_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_8_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_8_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_8_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_10_nl
      , while_and_132_nl , while_and_133_nl});
  assign while_or_11_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_11_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_9_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_136_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_11_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_137_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_9_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_9_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_9_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_11_nl
      , while_and_136_nl , while_and_137_nl});
  assign while_or_12_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_12_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_10_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_140_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_12_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_141_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_10_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_10_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_10_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_12_nl
      , while_and_140_nl , while_and_141_nl});
  assign while_or_13_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_13_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_11_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_144_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_13_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_145_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_11_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_11_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_11_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_13_nl
      , while_and_144_nl , while_and_145_nl});
  assign while_or_14_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_14_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_12_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_148_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_14_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_149_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_12_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_12_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_12_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_14_nl
      , while_and_148_nl , while_and_149_nl});
  assign while_or_15_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_15_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_13_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_152_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_15_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_153_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_13_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_13_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_13_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_15_nl
      , while_and_152_nl , while_and_153_nl});
  assign while_or_16_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_16_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_14_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_156_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_16_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_157_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_14_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_14_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_14_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_16_nl
      , while_and_156_nl , while_and_157_nl});
  assign while_or_17_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_17_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_15_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_160_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_17_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_161_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_15_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_15_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_15_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_17_nl
      , while_and_160_nl , while_and_161_nl});
  assign while_or_18_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_18_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_16_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_164_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_18_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_165_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_16_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_16_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_16_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_18_nl
      , while_and_164_nl , while_and_165_nl});
  assign while_or_19_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_19_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_17_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_168_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_19_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_169_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_17_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_17_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_17_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_19_nl
      , while_and_168_nl , while_and_169_nl});
  assign while_or_20_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_20_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_18_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_172_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_20_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_173_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_18_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_18_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_18_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_20_nl
      , while_and_172_nl , while_and_173_nl});
  assign while_or_21_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_21_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_19_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_176_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_21_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_177_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_19_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_19_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_19_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_21_nl
      , while_and_176_nl , while_and_177_nl});
  assign while_or_22_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_22_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_20_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_180_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_22_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_181_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_20_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_20_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_20_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_22_nl
      , while_and_180_nl , while_and_181_nl});
  assign while_or_23_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_23_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_21_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_184_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_23_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_185_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_21_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_21_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_21_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_23_nl
      , while_and_184_nl , while_and_185_nl});
  assign while_or_24_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_24_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_22_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_188_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_24_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_189_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_22_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_22_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_22_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_24_nl
      , while_and_188_nl , while_and_189_nl});
  assign while_or_25_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_25_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_23_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_192_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_25_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_193_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_23_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_23_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_23_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_25_nl
      , while_and_192_nl , while_and_193_nl});
  assign while_or_26_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_26_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_24_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_196_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_26_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_197_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_24_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_24_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_24_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_26_nl
      , while_and_196_nl , while_and_197_nl});
  assign while_or_27_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_27_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_25_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_200_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_27_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_201_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_25_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_25_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_25_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_27_nl
      , while_and_200_nl , while_and_201_nl});
  assign while_or_28_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_28_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_26_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_204_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_28_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_205_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_26_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_26_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_26_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_28_nl
      , while_and_204_nl , while_and_205_nl});
  assign while_or_29_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_29_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_27_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_208_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_29_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_209_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_27_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_27_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_27_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_29_nl
      , while_and_208_nl , while_and_209_nl});
  assign while_or_30_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_30_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_28_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_212_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_30_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_213_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_28_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_28_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_28_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_30_nl
      , while_and_212_nl , while_and_213_nl});
  assign while_or_31_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_31_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_29_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_216_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_31_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_217_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_29_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_29_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_29_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_31_nl
      , while_and_216_nl , while_and_217_nl});
  assign while_or_32_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_32_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_30_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_220_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_32_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_221_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_30_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_30_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_30_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_32_nl
      , while_and_220_nl , while_and_221_nl});
  assign while_or_33_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_33_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_31_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_224_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_33_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_225_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_31_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_31_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_31_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_33_nl
      , while_and_224_nl , while_and_225_nl});
  assign while_or_34_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_34_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_32_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_228_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_34_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_229_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_32_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_32_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_32_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_34_nl
      , while_and_228_nl , while_and_229_nl});
  assign while_or_35_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_35_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_33_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_232_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_35_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_233_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_33_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_33_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_33_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_35_nl
      , while_and_232_nl , while_and_233_nl});
  assign while_or_36_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_36_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_34_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_236_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_36_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_237_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_34_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_34_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_34_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_36_nl
      , while_and_236_nl , while_and_237_nl});
  assign while_or_37_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_37_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_35_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_240_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_37_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_241_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_35_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_35_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_35_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_37_nl
      , while_and_240_nl , while_and_241_nl});
  assign while_or_38_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_38_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_36_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_244_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_38_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_245_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_36_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_36_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_36_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_38_nl
      , while_and_244_nl , while_and_245_nl});
  assign while_or_39_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_39_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_37_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_248_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_39_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_249_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_37_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_37_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_37_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_39_nl
      , while_and_248_nl , while_and_249_nl});
  assign while_or_40_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_40_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_38_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_252_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_40_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_253_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_38_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_38_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_38_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_40_nl
      , while_and_252_nl , while_and_253_nl});
  assign while_or_41_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_41_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_39_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_256_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_41_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_257_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_39_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_39_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_39_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_41_nl
      , while_and_256_nl , while_and_257_nl});
  assign while_or_42_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_42_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_40_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_260_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_42_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_261_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_40_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_40_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_40_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_42_nl
      , while_and_260_nl , while_and_261_nl});
  assign while_or_43_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_43_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_41_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_264_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_43_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_265_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_41_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_41_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_41_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_43_nl
      , while_and_264_nl , while_and_265_nl});
  assign while_or_44_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_44_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_42_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_268_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_44_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_269_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_42_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_42_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_42_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_44_nl
      , while_and_268_nl , while_and_269_nl});
  assign while_or_45_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_45_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_43_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_272_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_45_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_273_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_43_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_43_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_43_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_45_nl
      , while_and_272_nl , while_and_273_nl});
  assign while_or_46_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_46_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_44_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_276_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_46_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_277_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_44_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_44_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_44_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_46_nl
      , while_and_276_nl , while_and_277_nl});
  assign while_or_47_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_47_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_45_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_280_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_47_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_281_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_45_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_45_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_45_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_47_nl
      , while_and_280_nl , while_and_281_nl});
  assign while_or_48_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_48_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_46_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_284_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_48_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_285_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_46_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_46_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_46_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_48_nl
      , while_and_284_nl , while_and_285_nl});
  assign while_or_49_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_49_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_47_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_288_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_49_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_289_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_47_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_47_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_47_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_49_nl
      , while_and_288_nl , while_and_289_nl});
  assign while_or_50_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_50_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_48_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_292_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_50_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_293_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_48_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_48_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_48_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_50_nl
      , while_and_292_nl , while_and_293_nl});
  assign while_or_51_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_51_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_49_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_296_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_51_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_297_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_49_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_49_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_49_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_51_nl
      , while_and_296_nl , while_and_297_nl});
  assign while_or_52_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_52_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_50_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_300_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_52_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_301_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_50_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_50_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_50_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_52_nl
      , while_and_300_nl , while_and_301_nl});
  assign while_or_53_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_53_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_51_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_304_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_53_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_305_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_51_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_51_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_51_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_53_nl
      , while_and_304_nl , while_and_305_nl});
  assign while_or_54_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_54_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_52_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_308_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_54_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_309_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_52_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_52_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_52_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_54_nl
      , while_and_308_nl , while_and_309_nl});
  assign while_or_55_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_55_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_53_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_312_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_55_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_313_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_53_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_53_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_53_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_55_nl
      , while_and_312_nl , while_and_313_nl});
  assign while_or_56_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_56_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_54_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_316_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_56_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_317_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_54_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_54_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_54_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_56_nl
      , while_and_316_nl , while_and_317_nl});
  assign while_or_57_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_57_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_55_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_320_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_57_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_321_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_55_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_55_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_55_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_57_nl
      , while_and_320_nl , while_and_321_nl});
  assign while_or_58_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_58_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_56_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_324_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_58_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_325_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_56_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_56_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_56_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_58_nl
      , while_and_324_nl , while_and_325_nl});
  assign while_or_59_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_59_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_57_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_328_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_59_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_329_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_57_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_57_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_57_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_59_nl
      , while_and_328_nl , while_and_329_nl});
  assign while_or_60_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_60_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_58_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_332_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_60_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_333_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_58_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_58_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_58_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_60_nl
      , while_and_332_nl , while_and_333_nl});
  assign while_or_61_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_61_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_59_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_336_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_61_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_337_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_59_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_59_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_59_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_61_nl
      , while_and_336_nl , while_and_337_nl});
  assign while_or_62_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_62_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_60_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_340_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_62_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_341_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_60_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_60_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_60_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_62_nl
      , while_and_340_nl , while_and_341_nl});
  assign while_or_63_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_63_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_61_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_344_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_63_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_345_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_61_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_61_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_61_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_63_nl
      , while_and_344_nl , while_and_345_nl});
  assign while_or_64_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_64_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_62_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_348_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_64_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_349_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_62_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_62_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_62_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_64_nl
      , while_and_348_nl , while_and_349_nl});
  assign while_or_65_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_65_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_63_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_352_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_65_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_353_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_63_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_63_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_63_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_65_nl
      , while_and_352_nl , while_and_353_nl});
  assign while_or_66_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_66_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_64_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_356_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_66_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_357_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_64_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_64_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_64_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_66_nl
      , while_and_356_nl , while_and_357_nl});
  assign while_or_67_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_67_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_65_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_360_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_67_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_361_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_65_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_65_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_65_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_67_nl
      , while_and_360_nl , while_and_361_nl});
  assign while_or_68_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_68_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_66_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_364_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_68_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_365_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_66_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_66_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_66_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_68_nl
      , while_and_364_nl , while_and_365_nl});
  assign while_or_69_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_69_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_67_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_368_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_69_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_369_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_67_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_67_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_67_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_69_nl
      , while_and_368_nl , while_and_369_nl});
  assign while_or_70_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_70_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_68_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_372_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_70_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_373_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_68_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_68_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_68_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_70_nl
      , while_and_372_nl , while_and_373_nl});
  assign while_or_71_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_71_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_69_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_376_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_71_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_377_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_69_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_69_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_69_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_71_nl
      , while_and_376_nl , while_and_377_nl});
  assign while_or_72_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_72_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_70_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_380_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_72_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_381_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_70_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_70_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_70_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_72_nl
      , while_and_380_nl , while_and_381_nl});
  assign while_or_73_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_73_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_71_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_384_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_73_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_385_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_71_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_71_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_71_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_73_nl
      , while_and_384_nl , while_and_385_nl});
  assign while_or_74_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_74_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_72_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_388_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_74_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_389_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_72_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_72_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_72_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_74_nl
      , while_and_388_nl , while_and_389_nl});
  assign while_or_75_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_75_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_73_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_392_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_75_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_393_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_73_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_73_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_73_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_75_nl
      , while_and_392_nl , while_and_393_nl});
  assign while_or_76_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_76_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_74_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_396_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_76_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_397_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_74_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_74_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_74_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_76_nl
      , while_and_396_nl , while_and_397_nl});
  assign while_or_77_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_77_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_75_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_400_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_77_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_401_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_75_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_75_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_75_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_77_nl
      , while_and_400_nl , while_and_401_nl});
  assign while_or_78_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_78_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_76_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_404_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_78_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_405_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_76_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_76_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_76_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_78_nl
      , while_and_404_nl , while_and_405_nl});
  assign while_or_79_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_79_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_77_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_408_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_79_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_409_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_77_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_77_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_77_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_79_nl
      , while_and_408_nl , while_and_409_nl});
  assign while_or_80_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_80_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_78_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_412_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_80_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_413_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_78_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_78_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_78_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_80_nl
      , while_and_412_nl , while_and_413_nl});
  assign while_or_81_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_81_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_79_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_416_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_81_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_417_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_79_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_79_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_79_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_81_nl
      , while_and_416_nl , while_and_417_nl});
  assign while_or_82_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_82_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_80_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_420_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_82_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_421_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_80_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_80_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_80_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_82_nl
      , while_and_420_nl , while_and_421_nl});
  assign while_or_83_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_83_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_81_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_424_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_83_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_425_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_81_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_81_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_81_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_83_nl
      , while_and_424_nl , while_and_425_nl});
  assign while_or_84_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_84_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_82_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_428_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_84_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_429_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_82_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_82_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_82_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_84_nl
      , while_and_428_nl , while_and_429_nl});
  assign while_or_85_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_85_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_83_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_432_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_85_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_433_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_83_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_83_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_83_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_85_nl
      , while_and_432_nl , while_and_433_nl});
  assign while_or_86_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_86_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_84_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_436_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_86_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_437_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_84_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_84_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_84_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_86_nl
      , while_and_436_nl , while_and_437_nl});
  assign while_or_87_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_87_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_85_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_440_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_87_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_441_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_85_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_85_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_85_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_87_nl
      , while_and_440_nl , while_and_441_nl});
  assign while_or_88_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_88_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_86_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_444_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_88_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_445_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_86_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_86_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_86_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_88_nl
      , while_and_444_nl , while_and_445_nl});
  assign while_or_89_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_89_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_87_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_448_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_89_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_449_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_87_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_87_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_87_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_89_nl
      , while_and_448_nl , while_and_449_nl});
  assign while_or_90_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_90_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_88_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_452_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_90_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_453_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_88_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_88_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_88_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_90_nl
      , while_and_452_nl , while_and_453_nl});
  assign while_or_91_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_91_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_89_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_456_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_91_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_457_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_89_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_89_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_89_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_91_nl
      , while_and_456_nl , while_and_457_nl});
  assign while_or_92_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_92_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_90_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_460_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_92_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_461_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_90_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_90_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_90_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_92_nl
      , while_and_460_nl , while_and_461_nl});
  assign while_or_93_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_93_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_91_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_464_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_93_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_465_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_91_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_91_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_91_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_93_nl
      , while_and_464_nl , while_and_465_nl});
  assign while_or_94_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_94_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_92_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_468_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_94_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_469_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_92_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_92_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_92_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_94_nl
      , while_and_468_nl , while_and_469_nl});
  assign while_or_95_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_95_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_93_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_472_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_95_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_473_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_93_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_93_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_93_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_95_nl
      , while_and_472_nl , while_and_473_nl});
  assign while_or_96_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_96_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_94_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_476_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_96_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_477_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_94_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_94_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_94_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_96_nl
      , while_and_476_nl , while_and_477_nl});
  assign while_or_97_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_97_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_95_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_480_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_97_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_481_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_95_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_95_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_95_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_97_nl
      , while_and_480_nl , while_and_481_nl});
  assign while_or_98_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_98_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_96_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_484_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_98_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_485_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_96_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_96_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_96_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_98_nl
      , while_and_484_nl , while_and_485_nl});
  assign while_or_99_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_99_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_97_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_488_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_99_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_489_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_97_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_97_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_97_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_99_nl
      , while_and_488_nl , while_and_489_nl});
  assign while_or_100_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_100_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_98_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_492_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_100_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_493_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_98_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_98_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_98_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_100_nl
      , while_and_492_nl , while_and_493_nl});
  assign while_or_101_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_101_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_99_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_496_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_101_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_497_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_99_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_99_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_99_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_101_nl
      , while_and_496_nl , while_and_497_nl});
  assign while_or_102_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_102_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_100_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_500_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_102_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_501_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_100_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_100_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_100_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_102_nl
      , while_and_500_nl , while_and_501_nl});
  assign while_or_103_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_103_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_101_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_504_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_103_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_505_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_101_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_101_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_101_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_103_nl
      , while_and_504_nl , while_and_505_nl});
  assign while_or_104_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_104_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_102_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_508_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_104_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_509_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_102_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_102_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_102_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_104_nl
      , while_and_508_nl , while_and_509_nl});
  assign while_or_105_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_105_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_103_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_512_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_105_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_513_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_103_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_103_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_103_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_105_nl
      , while_and_512_nl , while_and_513_nl});
  assign while_or_106_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_106_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_104_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_516_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_106_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_517_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_104_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_104_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_104_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_106_nl
      , while_and_516_nl , while_and_517_nl});
  assign while_or_107_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_107_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_105_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_520_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_107_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_521_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_105_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_105_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_105_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_107_nl
      , while_and_520_nl , while_and_521_nl});
  assign while_or_108_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_108_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_106_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_524_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_108_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_525_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_106_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_106_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_106_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_108_nl
      , while_and_524_nl , while_and_525_nl});
  assign while_or_109_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_109_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_107_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_528_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_109_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_529_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_107_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_107_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_107_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_109_nl
      , while_and_528_nl , while_and_529_nl});
  assign while_or_110_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_110_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_108_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_532_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_110_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_533_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_108_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_108_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_108_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_110_nl
      , while_and_532_nl , while_and_533_nl});
  assign while_or_111_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_111_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_109_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_536_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_111_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_537_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_109_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_109_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_109_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_111_nl
      , while_and_536_nl , while_and_537_nl});
  assign while_or_112_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_112_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_110_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_540_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_112_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_541_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_110_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_110_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_110_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_112_nl
      , while_and_540_nl , while_and_541_nl});
  assign while_or_113_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_113_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_111_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_544_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_113_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_545_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_111_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_111_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_111_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_113_nl
      , while_and_544_nl , while_and_545_nl});
  assign while_or_114_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_114_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_112_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_548_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_114_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_549_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_112_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_112_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_112_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_114_nl
      , while_and_548_nl , while_and_549_nl});
  assign while_or_115_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_115_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_113_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_552_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_115_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_553_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_113_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_113_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_113_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_115_nl
      , while_and_552_nl , while_and_553_nl});
  assign while_or_116_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_116_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_114_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_556_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_116_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_557_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_114_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_114_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_114_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_116_nl
      , while_and_556_nl , while_and_557_nl});
  assign while_or_117_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_117_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_115_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_560_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_117_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_561_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_115_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_115_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_115_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_117_nl
      , while_and_560_nl , while_and_561_nl});
  assign while_or_118_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_118_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_116_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_564_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_118_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_565_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_116_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_116_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_116_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_118_nl
      , while_and_564_nl , while_and_565_nl});
  assign while_or_119_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_119_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_117_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_568_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_119_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_569_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_117_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_117_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_117_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_119_nl
      , while_and_568_nl , while_and_569_nl});
  assign while_or_120_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_120_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_118_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_572_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_120_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_573_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_118_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_118_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_118_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_120_nl
      , while_and_572_nl , while_and_573_nl});
  assign while_or_121_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_121_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_119_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_576_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_121_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_577_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_119_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_119_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_119_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_121_nl
      , while_and_576_nl , while_and_577_nl});
  assign while_or_122_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_122_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_120_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_580_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_122_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_581_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_120_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_120_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_120_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_122_nl
      , while_and_580_nl , while_and_581_nl});
  assign while_or_123_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_123_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_121_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_584_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_123_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_585_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_121_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_121_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_121_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_123_nl
      , while_and_584_nl , while_and_585_nl});
  assign while_or_124_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_124_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_122_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_588_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_124_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_589_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_122_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_122_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_122_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_124_nl
      , while_and_588_nl , while_and_589_nl});
  assign while_or_125_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_125_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_123_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_592_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_125_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_593_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_123_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_123_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_123_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_125_nl
      , while_and_592_nl , while_and_593_nl});
  assign while_or_126_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_126_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_124_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_596_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_126_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_597_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_124_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_124_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_124_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_126_nl
      , while_and_596_nl , while_and_597_nl});
  assign while_or_127_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_127_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_125_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_600_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_127_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_601_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_125_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_125_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_125_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_127_nl
      , while_and_600_nl , while_and_601_nl});
  assign while_or_128_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_128_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_126_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_604_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_128_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_605_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_126_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_126_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_126_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_128_nl
      , while_and_604_nl , while_and_605_nl});
  assign while_or_129_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_129_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_127_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_608_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_129_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_609_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_127_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_127_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_127_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_129_nl
      , while_and_608_nl , while_and_609_nl});
  assign while_or_130_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_130_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_128_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_612_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_130_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_613_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_128_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_128_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_128_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_130_nl
      , while_and_612_nl , while_and_613_nl});
  assign while_or_131_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_131_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_129_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_616_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_131_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_617_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_129_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_129_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_129_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_131_nl
      , while_and_616_nl , while_and_617_nl});
  assign while_or_132_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_132_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_130_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_620_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_132_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_621_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_130_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_130_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_130_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_132_nl
      , while_and_620_nl , while_and_621_nl});
  assign while_or_133_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_133_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_131_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_624_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_133_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_625_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_131_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_131_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_131_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_133_nl
      , while_and_624_nl , while_and_625_nl});
  assign while_or_134_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_134_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_132_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_628_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_134_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_629_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_132_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_132_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_132_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_134_nl
      , while_and_628_nl , while_and_629_nl});
  assign while_or_135_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_135_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_133_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_632_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_135_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_633_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_133_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_133_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_133_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_135_nl
      , while_and_632_nl , while_and_633_nl});
  assign while_or_136_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_136_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_134_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_636_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_136_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_637_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_134_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_134_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_134_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_136_nl
      , while_and_636_nl , while_and_637_nl});
  assign while_or_137_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_137_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_135_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_640_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_137_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_641_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_135_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_135_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_135_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_137_nl
      , while_and_640_nl , while_and_641_nl});
  assign while_or_138_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_138_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_136_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_644_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_138_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_645_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_136_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_136_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_136_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_138_nl
      , while_and_644_nl , while_and_645_nl});
  assign while_or_139_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_139_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_137_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_648_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_139_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_649_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_137_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_137_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_137_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_139_nl
      , while_and_648_nl , while_and_649_nl});
  assign while_or_140_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_140_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_138_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_652_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_140_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_653_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_138_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_138_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_138_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_140_nl
      , while_and_652_nl , while_and_653_nl});
  assign while_or_141_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_141_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_139_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_656_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_141_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_657_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_139_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_139_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_139_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_141_nl
      , while_and_656_nl , while_and_657_nl});
  assign while_or_142_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_142_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_140_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_660_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_142_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_661_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_140_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_140_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_140_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_142_nl
      , while_and_660_nl , while_and_661_nl});
  assign while_or_143_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_143_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_141_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_664_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_143_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_665_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_141_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_141_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_141_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_143_nl
      , while_and_664_nl , while_and_665_nl});
  assign while_or_144_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_144_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_142_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_668_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_144_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_669_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_142_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_142_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_142_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_144_nl
      , while_and_668_nl , while_and_669_nl});
  assign while_or_145_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_145_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_143_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_672_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_145_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_673_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_143_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_143_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_143_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_145_nl
      , while_and_672_nl , while_and_673_nl});
  assign while_or_146_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_146_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_144_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_676_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_146_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_677_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_144_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_144_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_144_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_146_nl
      , while_and_676_nl , while_and_677_nl});
  assign while_or_147_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_147_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_145_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_680_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_147_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_681_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_145_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_145_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_145_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_147_nl
      , while_and_680_nl , while_and_681_nl});
  assign while_or_148_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_148_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_146_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_684_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_148_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_685_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_146_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_146_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_146_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_148_nl
      , while_and_684_nl , while_and_685_nl});
  assign while_or_149_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_149_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_147_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_688_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_149_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_689_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_147_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_147_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_147_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_149_nl
      , while_and_688_nl , while_and_689_nl});
  assign while_or_150_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_150_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_148_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_692_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_150_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_693_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_148_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_148_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_148_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_150_nl
      , while_and_692_nl , while_and_693_nl});
  assign while_or_151_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_151_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_149_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_696_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_151_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_697_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_149_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_149_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_149_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_151_nl
      , while_and_696_nl , while_and_697_nl});
  assign while_or_152_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_152_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_150_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_700_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_152_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_701_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_150_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_150_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_150_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_152_nl
      , while_and_700_nl , while_and_701_nl});
  assign while_or_153_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_153_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_151_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_704_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_153_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_705_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_151_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_151_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_151_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_153_nl
      , while_and_704_nl , while_and_705_nl});
  assign while_or_154_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_154_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_152_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_708_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_154_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_709_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_152_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_152_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_152_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_154_nl
      , while_and_708_nl , while_and_709_nl});
  assign while_or_155_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_155_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_153_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_712_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_155_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_713_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_153_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_153_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_153_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_155_nl
      , while_and_712_nl , while_and_713_nl});
  assign while_or_156_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_156_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_154_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_716_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_156_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_717_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_154_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_154_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_154_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_156_nl
      , while_and_716_nl , while_and_717_nl});
  assign while_or_157_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_157_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_155_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_720_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_157_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_721_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_155_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_155_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_155_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_157_nl
      , while_and_720_nl , while_and_721_nl});
  assign while_or_158_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_158_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_156_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_724_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_158_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_725_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_156_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_156_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_156_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_158_nl
      , while_and_724_nl , while_and_725_nl});
  assign while_or_159_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_159_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_157_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_728_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_159_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_729_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_157_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_157_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_157_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_159_nl
      , while_and_728_nl , while_and_729_nl});
  assign while_or_160_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_160_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_158_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_732_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_160_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_733_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_158_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_158_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_158_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_160_nl
      , while_and_732_nl , while_and_733_nl});
  assign while_or_161_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_161_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_159_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_736_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_161_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_737_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_159_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_159_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_159_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_161_nl
      , while_and_736_nl , while_and_737_nl});
  assign while_or_162_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_162_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_160_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_740_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_162_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_741_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_160_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_160_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_160_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_162_nl
      , while_and_740_nl , while_and_741_nl});
  assign while_or_163_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_163_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_161_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_744_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_163_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_745_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_161_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_161_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_161_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_163_nl
      , while_and_744_nl , while_and_745_nl});
  assign while_or_164_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_164_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_162_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_748_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_164_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_749_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_162_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_162_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_162_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_164_nl
      , while_and_748_nl , while_and_749_nl});
  assign while_or_165_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_165_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_163_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_752_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_165_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_753_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_163_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_163_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_163_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_165_nl
      , while_and_752_nl , while_and_753_nl});
  assign while_or_166_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_166_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_164_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_756_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_166_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_757_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_164_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_164_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_164_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_166_nl
      , while_and_756_nl , while_and_757_nl});
  assign while_or_167_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_167_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_165_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_760_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_167_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_761_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_165_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_165_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_165_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_167_nl
      , while_and_760_nl , while_and_761_nl});
  assign while_or_168_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_168_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_166_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_764_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_168_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_765_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_166_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_166_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_166_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_168_nl
      , while_and_764_nl , while_and_765_nl});
  assign while_or_169_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_169_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_167_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_768_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_169_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_769_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_167_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_167_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_167_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_169_nl
      , while_and_768_nl , while_and_769_nl});
  assign while_or_170_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_170_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_168_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_772_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_170_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_773_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_168_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_168_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_168_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_170_nl
      , while_and_772_nl , while_and_773_nl});
  assign while_or_171_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_171_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_169_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_776_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_171_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_777_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_169_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_169_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_169_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_171_nl
      , while_and_776_nl , while_and_777_nl});
  assign while_or_172_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_172_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_170_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_780_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_172_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_781_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_170_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_170_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_170_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_172_nl
      , while_and_780_nl , while_and_781_nl});
  assign while_or_173_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_173_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_171_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_784_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_173_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_785_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_171_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_171_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_171_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_173_nl
      , while_and_784_nl , while_and_785_nl});
  assign while_or_174_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_174_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_172_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_788_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_174_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_789_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_172_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_172_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_172_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_174_nl
      , while_and_788_nl , while_and_789_nl});
  assign while_or_175_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_175_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_173_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_792_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_175_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_793_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_173_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_173_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_173_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_175_nl
      , while_and_792_nl , while_and_793_nl});
  assign while_or_176_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_176_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_174_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_796_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_176_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_797_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_174_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_174_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_174_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_176_nl
      , while_and_796_nl , while_and_797_nl});
  assign while_or_177_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_177_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_175_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_800_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_177_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_801_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_175_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_175_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_175_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_177_nl
      , while_and_800_nl , while_and_801_nl});
  assign while_or_178_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_178_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_176_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_804_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_178_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_805_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_176_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_176_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_176_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_178_nl
      , while_and_804_nl , while_and_805_nl});
  assign while_or_179_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_179_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_177_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_808_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_179_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_809_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_177_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_177_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_177_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_179_nl
      , while_and_808_nl , while_and_809_nl});
  assign while_or_180_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_180_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_178_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_812_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_180_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_813_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_178_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_178_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_178_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_180_nl
      , while_and_812_nl , while_and_813_nl});
  assign while_or_181_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_181_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_179_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_816_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_181_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_817_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_179_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_179_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_179_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_181_nl
      , while_and_816_nl , while_and_817_nl});
  assign while_or_182_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_182_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_180_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_820_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_182_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_821_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_180_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_180_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_180_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_182_nl
      , while_and_820_nl , while_and_821_nl});
  assign while_or_183_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_183_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_181_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_824_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_183_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_825_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_181_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_181_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_181_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_183_nl
      , while_and_824_nl , while_and_825_nl});
  assign while_or_184_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_184_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_182_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_828_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_184_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_829_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_182_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_182_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_182_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_184_nl
      , while_and_828_nl , while_and_829_nl});
  assign while_or_185_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_185_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_183_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_832_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_185_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_833_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_183_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_183_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_183_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_185_nl
      , while_and_832_nl , while_and_833_nl});
  assign while_or_186_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_186_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_184_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_836_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_186_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_837_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_184_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_184_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_184_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_186_nl
      , while_and_836_nl , while_and_837_nl});
  assign while_or_187_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_187_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_185_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_840_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_187_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_841_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_185_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_185_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_185_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_187_nl
      , while_and_840_nl , while_and_841_nl});
  assign while_or_188_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_188_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_186_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_844_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_188_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_845_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_186_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_186_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_186_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_188_nl
      , while_and_844_nl , while_and_845_nl});
  assign while_or_189_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_189_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_187_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_848_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_189_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_849_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_187_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_187_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_187_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_189_nl
      , while_and_848_nl , while_and_849_nl});
  assign while_or_190_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_190_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_188_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_852_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_190_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_853_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_188_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_188_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_188_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_190_nl
      , while_and_852_nl , while_and_853_nl});
  assign while_or_191_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_191_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_189_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_856_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_191_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_857_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_189_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_189_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_189_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_191_nl
      , while_and_856_nl , while_and_857_nl});
  assign while_or_192_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_192_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_190_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_860_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_192_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_861_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_190_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_190_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_190_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_192_nl
      , while_and_860_nl , while_and_861_nl});
  assign while_or_193_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_193_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_191_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_864_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_193_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_865_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_191_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_191_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_191_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_193_nl
      , while_and_864_nl , while_and_865_nl});
  assign while_or_194_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_194_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_192_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_868_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_194_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_869_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_192_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_192_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_192_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_194_nl
      , while_and_868_nl , while_and_869_nl});
  assign while_or_195_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_195_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_193_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_872_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_195_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_873_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_193_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_193_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_193_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_195_nl
      , while_and_872_nl , while_and_873_nl});
  assign while_or_196_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_196_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_194_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_876_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_196_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_877_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_194_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_194_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_194_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_196_nl
      , while_and_876_nl , while_and_877_nl});
  assign while_or_197_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_197_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_195_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_880_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_197_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_881_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_195_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_195_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_195_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_197_nl
      , while_and_880_nl , while_and_881_nl});
  assign while_or_198_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_198_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_196_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_884_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_198_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_885_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_196_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_196_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_196_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_198_nl
      , while_and_884_nl , while_and_885_nl});
  assign while_or_199_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_199_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_197_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_888_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_199_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_889_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_197_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_197_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_197_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_199_nl
      , while_and_888_nl , while_and_889_nl});
  assign while_or_200_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_200_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_198_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_892_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_200_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_893_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_198_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_198_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_198_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_200_nl
      , while_and_892_nl , while_and_893_nl});
  assign while_or_201_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_201_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_199_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_896_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_201_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_897_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_199_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_199_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_199_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_201_nl
      , while_and_896_nl , while_and_897_nl});
  assign while_or_202_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_202_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_200_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_900_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_202_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_901_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_200_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_200_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_200_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_202_nl
      , while_and_900_nl , while_and_901_nl});
  assign while_or_203_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_203_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_201_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_904_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_203_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_905_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_201_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_201_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_201_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_203_nl
      , while_and_904_nl , while_and_905_nl});
  assign while_or_204_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_204_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_202_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_908_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_204_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_909_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_202_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_202_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_202_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_204_nl
      , while_and_908_nl , while_and_909_nl});
  assign while_or_205_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_205_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_203_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_912_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_205_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_913_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_203_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_203_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_203_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_205_nl
      , while_and_912_nl , while_and_913_nl});
  assign while_or_206_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_206_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_204_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_916_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_206_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_917_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_204_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_204_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_204_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_206_nl
      , while_and_916_nl , while_and_917_nl});
  assign while_or_207_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_207_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_205_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_920_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_207_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_921_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_205_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_205_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_205_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_207_nl
      , while_and_920_nl , while_and_921_nl});
  assign while_or_208_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_208_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_206_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_924_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_208_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_925_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_206_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_206_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_206_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_208_nl
      , while_and_924_nl , while_and_925_nl});
  assign while_or_209_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_209_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_207_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_928_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_209_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_929_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_207_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_207_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_207_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_209_nl
      , while_and_928_nl , while_and_929_nl});
  assign while_or_210_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_210_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_208_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_932_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_210_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_933_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_208_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_208_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_208_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_210_nl
      , while_and_932_nl , while_and_933_nl});
  assign while_or_211_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_211_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_209_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_936_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_211_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_937_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_209_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_209_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_209_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_211_nl
      , while_and_936_nl , while_and_937_nl});
  assign while_or_212_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_212_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_210_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_940_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_212_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_941_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_210_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_210_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_210_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_212_nl
      , while_and_940_nl , while_and_941_nl});
  assign while_or_213_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_213_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_211_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_944_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_213_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_945_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_211_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_211_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_211_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_213_nl
      , while_and_944_nl , while_and_945_nl});
  assign while_or_214_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_214_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_212_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_948_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_214_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_949_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_212_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_212_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_212_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_214_nl
      , while_and_948_nl , while_and_949_nl});
  assign while_or_215_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_215_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_213_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_952_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_215_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_953_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_213_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_213_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_213_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_215_nl
      , while_and_952_nl , while_and_953_nl});
  assign while_or_216_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_216_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_214_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_956_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_216_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_957_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_214_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_214_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_214_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_216_nl
      , while_and_956_nl , while_and_957_nl});
  assign while_or_217_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_217_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_215_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_960_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_217_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_961_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_215_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_215_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_215_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_217_nl
      , while_and_960_nl , while_and_961_nl});
  assign while_or_218_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_218_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_216_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_964_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_218_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_965_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_216_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_216_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_216_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_218_nl
      , while_and_964_nl , while_and_965_nl});
  assign while_or_219_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_219_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_217_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_968_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_219_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_969_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_217_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_217_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_217_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_219_nl
      , while_and_968_nl , while_and_969_nl});
  assign while_or_220_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_220_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_218_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_972_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_220_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_973_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_218_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_218_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_218_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_220_nl
      , while_and_972_nl , while_and_973_nl});
  assign while_or_221_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_221_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_219_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_976_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_221_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_977_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_219_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_219_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_219_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_221_nl
      , while_and_976_nl , while_and_977_nl});
  assign while_or_222_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_222_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_220_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_980_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_222_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_981_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_220_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_220_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_220_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_222_nl
      , while_and_980_nl , while_and_981_nl});
  assign while_or_223_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_223_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_221_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_984_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_223_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_985_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_221_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_221_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_221_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_223_nl
      , while_and_984_nl , while_and_985_nl});
  assign while_or_224_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_224_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_222_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_988_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_224_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_989_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_222_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_222_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_222_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_224_nl
      , while_and_988_nl , while_and_989_nl});
  assign while_or_225_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_225_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_223_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_992_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_225_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_993_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_223_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_223_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_223_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_225_nl
      , while_and_992_nl , while_and_993_nl});
  assign while_or_226_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_226_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_224_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_996_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_226_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_997_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_224_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_224_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_224_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_226_nl
      , while_and_996_nl , while_and_997_nl});
  assign while_or_227_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_227_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_225_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1000_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_227_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1001_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_225_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_225_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_225_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_227_nl
      , while_and_1000_nl , while_and_1001_nl});
  assign while_or_228_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_228_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_226_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1004_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_228_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1005_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_226_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_226_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_226_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_228_nl
      , while_and_1004_nl , while_and_1005_nl});
  assign while_or_229_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_229_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_227_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1008_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_229_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1009_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_227_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_227_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_227_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_229_nl
      , while_and_1008_nl , while_and_1009_nl});
  assign while_or_230_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_230_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_228_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1012_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_230_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1013_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_228_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_228_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_228_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_230_nl
      , while_and_1012_nl , while_and_1013_nl});
  assign while_or_231_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_231_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_229_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1016_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_231_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1017_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_229_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_229_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_229_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_231_nl
      , while_and_1016_nl , while_and_1017_nl});
  assign while_or_232_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_232_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_230_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1020_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_232_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1021_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_230_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_230_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_230_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_232_nl
      , while_and_1020_nl , while_and_1021_nl});
  assign while_or_233_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_233_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_231_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1024_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_233_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1025_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_231_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_231_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_231_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_233_nl
      , while_and_1024_nl , while_and_1025_nl});
  assign while_or_234_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_234_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_232_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1028_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_234_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1029_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_232_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_232_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_232_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_234_nl
      , while_and_1028_nl , while_and_1029_nl});
  assign while_or_235_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_235_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_233_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1032_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_235_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1033_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_233_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_233_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_233_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_235_nl
      , while_and_1032_nl , while_and_1033_nl});
  assign while_or_236_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_236_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_234_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1036_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_236_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1037_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_234_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_234_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_234_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_236_nl
      , while_and_1036_nl , while_and_1037_nl});
  assign while_or_237_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_237_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_235_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1040_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_237_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1041_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_235_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_235_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_235_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_237_nl
      , while_and_1040_nl , while_and_1041_nl});
  assign while_or_238_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_238_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_236_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1044_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_238_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1045_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_236_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_236_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_236_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_238_nl
      , while_and_1044_nl , while_and_1045_nl});
  assign while_or_239_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_239_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_237_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1048_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_239_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1049_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_237_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_237_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_237_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_239_nl
      , while_and_1048_nl , while_and_1049_nl});
  assign while_or_240_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_240_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_238_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1052_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_240_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1053_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_238_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_238_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_238_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_240_nl
      , while_and_1052_nl , while_and_1053_nl});
  assign while_or_241_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_241_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_239_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1056_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_241_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1057_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_239_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_239_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_239_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_241_nl
      , while_and_1056_nl , while_and_1057_nl});
  assign while_or_242_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_242_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_240_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1060_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_242_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1061_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_240_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_240_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_240_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_242_nl
      , while_and_1060_nl , while_and_1061_nl});
  assign while_or_243_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_243_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_241_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1064_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_243_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1065_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_241_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_241_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_241_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_243_nl
      , while_and_1064_nl , while_and_1065_nl});
  assign while_or_244_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_244_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_242_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1068_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_244_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1069_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_242_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_242_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_242_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_244_nl
      , while_and_1068_nl , while_and_1069_nl});
  assign while_or_245_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_245_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_243_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1072_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_245_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1073_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_243_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_243_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_243_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_245_nl
      , while_and_1072_nl , while_and_1073_nl});
  assign while_or_246_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_246_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_244_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1076_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_246_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1077_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_244_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_244_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_244_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_246_nl
      , while_and_1076_nl , while_and_1077_nl});
  assign while_or_247_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_247_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_245_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1080_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_247_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1081_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_245_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_245_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_245_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_247_nl
      , while_and_1080_nl , while_and_1081_nl});
  assign while_or_248_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_248_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_246_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1084_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_248_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1085_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_246_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_246_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_246_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_248_nl
      , while_and_1084_nl , while_and_1085_nl});
  assign while_or_249_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_249_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_247_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1088_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_249_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1089_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_247_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_247_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_247_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_249_nl
      , while_and_1088_nl , while_and_1089_nl});
  assign while_or_250_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_250_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_248_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1092_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_250_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1093_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_248_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_248_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_248_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_250_nl
      , while_and_1092_nl , while_and_1093_nl});
  assign while_or_251_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_251_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_249_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1096_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_251_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1097_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_249_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_249_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_249_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_251_nl
      , while_and_1096_nl , while_and_1097_nl});
  assign while_or_252_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_252_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_250_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1100_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_252_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1101_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_250_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_250_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_250_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_252_nl
      , while_and_1100_nl , while_and_1101_nl});
  assign while_or_253_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_253_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_251_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1104_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_253_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1105_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_251_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_251_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_251_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_253_nl
      , while_and_1104_nl , while_and_1105_nl});
  assign while_or_254_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_254_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_252_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1108_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_254_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1109_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_252_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_252_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_252_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_254_nl
      , while_and_1108_nl , while_and_1109_nl});
  assign while_or_255_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_255_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_253_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1112_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_255_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1113_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_253_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_253_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_253_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_255_nl
      , while_and_1112_nl , while_and_1113_nl});
  assign while_or_256_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_256_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_254_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1116_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_256_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1117_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_254_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_254_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_254_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_256_nl
      , while_and_1116_nl , while_and_1117_nl});
  assign while_or_257_nl = (~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_257_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_255_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1120_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_257_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign while_and_1121_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_255_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign input_mem_banks_bank_a_255_sva_dfm_2_mx0w0 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_255_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {while_or_257_nl
      , while_and_1120_nl , while_and_1121_nl});
  assign PECore_PushAxiRsp_mux_24_nl = MUX_s_1_2_2(reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse,
      PECore_PushAxiRsp_mux_10_itm_1, rva_in_reg_rw_sva_5);
  assign PECore_PushAxiRsp_if_else_mux_10_mx0w2 = MUX_s_1_2_2(PECore_PushAxiRsp_mux_24_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1);
  assign rva_out_reg_data_62_56_sva_dfm_6_mx1 = MUX_v_7_2_2(rva_out_reg_data_62_56_sva_dfm_4_1,
      rva_out_reg_data_62_56_sva_dfm_6, or_dcpl_283);
  assign rva_out_reg_data_35_32_sva_dfm_6_mx1 = MUX_v_4_2_2(rva_out_reg_data_35_32_sva_dfm_4_1,
      rva_out_reg_data_35_32_sva_dfm_6, or_dcpl_283);
  assign pe_manager_base_input_sva_mx1_7_0 = MUX_v_8_2_2((pe_manager_base_input_sva[7:0]),
      (pe_manager_base_input_sva_dfm_3_1[7:0]), while_stage_0_3);
  assign pe_manager_base_input_sva_mx2 = MUX_v_15_2_2(pe_manager_base_input_sva,
      pe_manager_base_input_sva_dfm_3_1, while_stage_0_3);
  assign PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
      & PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3
      | and_301_cse);
  assign PECore_RunScale_PECore_RunScale_if_and_1_svs_1 = (state_mux_1_cse[0]) &
      state_0_sva_mx1 & (~ (state_mux_1_cse[1]));
  assign PECore_DecodeAxiRead_switch_lp_nor_tmp_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_DecodeAxiRead_switch_lp_nor_9_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 | PECore_DecodeAxiRead_switch_lp_nor_tmp_10);
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1 = ~(input_read_req_valid_lpi_1_dfm_1_10
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_sva_1
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0 = MUX_v_64_2_2(weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0 = MUX_v_56_2_2(weight_mem_banks_read_1_read_data_lpi_1_dfm_1_63_8,
      (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63:8]), weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2});
  assign weight_mem_banks_load_store_1_for_else_else_and_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_or_nl = (weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1);
  assign weight_mem_banks_load_store_1_for_else_else_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9 = MUX1HOT_v_8_6_2(BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1,
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1,
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[7:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[7:0]),
      {weight_mem_banks_load_store_1_for_else_else_and_nl , weight_mem_banks_load_store_1_for_else_else_or_nl
      , weight_mem_banks_load_store_1_for_else_else_and_4_nl , weight_mem_banks_load_store_1_for_else_else_and_6_nl
      , weight_mem_banks_load_store_1_for_else_else_and_8_nl , weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {weight_mem_run_3_for_5_and_182_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_35_nl = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_000000
      = MUX_v_8_2_2(8'b00000000, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_35_nl,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_89_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_89_nl , weight_mem_run_3_for_5_asn_324
      , weight_mem_run_3_for_5_asn_326 , PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5
      , weight_mem_run_3_for_5_asn_328 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_2 , weight_mem_run_3_for_5_asn_330});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_81_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_81_nl , weight_mem_run_3_for_5_asn_324
      , weight_mem_run_3_for_5_asn_326 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1
      , weight_mem_run_3_for_5_asn_328 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_2
      , PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 , PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_73_cse = reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_73_cse , weight_mem_run_3_for_5_asn_324
      , weight_mem_run_3_for_5_asn_326 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_2
      , weight_mem_run_3_for_5_asn_328 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_73_cse , weight_mem_run_3_for_5_asn_324
      , weight_mem_run_3_for_5_asn_326 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2
      , weight_mem_run_3_for_5_asn_328 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2:1]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1 = (~(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_sva_1 | mux_160_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_sva_1 & (~ mux_160_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_2_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_sva_1) & not_tmp_425;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_sva_1 & not_tmp_425;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_sva_1) & and_dcpl_632;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_sva_1 & and_dcpl_632;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]),
      {mux_tmp_153 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_2_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_sva_1,
      {mux_tmp_153 , (~ mux_160_itm) , not_tmp_425 , and_dcpl_632});
  assign and_887_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  assign and_889_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  assign and_888_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  assign and_890_cse = weight_mem_read_arbxbar_arbiters_next_7_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign and_893_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) & while_mux_1303_tmp;
  assign and_892_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) & while_mux_1301_tmp;
  assign and_891_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) & while_mux_1304_tmp;
  assign and_894_cse = while_mux_1302_tmp & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign nor_419_nl = ~(and_887_cse | and_888_cse | and_889_cse | and_890_cse | or_tmp_209);
  assign nor_420_nl = ~(and_891_cse | and_892_cse | and_893_cse | and_894_cse | mux_tmp_152);
  assign mux_175_nl = MUX_s_1_2_2(nor_419_nl, nor_420_nl, while_stage_0_5);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl,
      mux_175_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 | mux_193_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 & (~ mux_193_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 | mux_207_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 & (~ mux_207_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1) & and_dcpl_634;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 & and_dcpl_634;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]),
      {mux_tmp_178 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1,
      {mux_tmp_178 , (~ mux_193_itm) , (~ mux_207_itm) , and_dcpl_634});
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  assign mux_216_nl = MUX_s_1_2_2(or_tmp_292, or_tmp_287, while_stage_0_5);
  assign or_581_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | or_tmp_292;
  assign or_576_nl = while_mux_1291_tmp | or_tmp_287;
  assign mux_215_nl = MUX_s_1_2_2(or_581_nl, or_576_nl, while_stage_0_5);
  assign mux_217_nl = MUX_s_1_2_2(mux_216_nl, mux_215_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl,
      mux_217_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 | mux_235_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 & (~ mux_235_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 | mux_244_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 & (~ mux_244_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1) & and_dcpl_637;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 & and_dcpl_637;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]),
      {mux_tmp_220 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1,
      {mux_tmp_220 , (~ mux_235_itm) , (~ mux_244_itm) , and_dcpl_637});
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl,
      mux_tmp_239);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1) & and_dcpl_642;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 & and_dcpl_642;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1) & and_dcpl_643;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 & and_dcpl_643;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1) & and_dcpl_644;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 & and_dcpl_644;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]),
      {and_dcpl_639 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_18_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_20_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1,
      {and_dcpl_639 , and_dcpl_642 , and_dcpl_643 , and_dcpl_644});
  assign operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 | mux_264_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 & (~ mux_264_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 | mux_277_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 & (~ mux_277_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1) & and_dcpl_647;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 & and_dcpl_647;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]),
      {mux_tmp_255 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1,
      {mux_tmp_255 , (~ mux_264_itm) , (~ mux_277_itm) , and_dcpl_647});
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_4_sva_1;
  assign mux_286_nl = MUX_s_1_2_2(or_tmp_373, or_tmp_368, while_stage_0_5);
  assign or_665_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1
      | or_tmp_373;
  assign or_660_nl = while_mux_1270_tmp | or_tmp_368;
  assign mux_285_nl = MUX_s_1_2_2(or_665_nl, or_660_nl, while_stage_0_5);
  assign mux_287_nl = MUX_s_1_2_2(mux_286_nl, mux_285_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl,
      mux_287_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_3_nl
      = weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 | mux_295_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 & (~ mux_295_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_32_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1) & and_dcpl_648;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 & and_dcpl_648;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1) & and_dcpl_652;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 & and_dcpl_652;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_3_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]),
      {mux_tmp_290 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_32_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1,
      {mux_tmp_290 , (~ mux_295_itm) , and_dcpl_648 , and_dcpl_652});
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign mux_304_nl = MUX_s_1_2_2(mux_tmp_297, mux_tmp_296, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign nor_421_nl = ~(mux_304_nl | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl,
      nor_421_nl);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      = weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | (weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]));
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_41_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_111_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_103_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_99_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_79_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_75_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_67_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_63_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_55_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_51_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_43_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_39_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = (pe_manager_base_weight_sva_mx2[14:4])
      + PEManager_15U_GetWeightAddr_else_acc_3_1;
  assign PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1[10:0];
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1) & and_dcpl_655;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 & and_dcpl_655;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1) & and_dcpl_656;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 & and_dcpl_656;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1) & and_dcpl_657;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 & and_dcpl_657;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]),
      {weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_tmp
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_36_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_38_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1,
      {weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_tmp
      , and_dcpl_655 , and_dcpl_656 , and_dcpl_657});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_tmp,
      weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_tmp,
      weight_mem_read_arbxbar_xbar_1_for_3_2_operator_7_false_1_operator_7_false_1_or_tmp);
  assign operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_tmp
      = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_tmp
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_7_false_1_operator_7_false_1_or_tmp
      = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]));
  assign nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_4_mux_2_mx0w2
      = MUX_s_1_2_2((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]),
      operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1);
  assign nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_5_mux_2_mx0w3
      = MUX_s_1_2_2((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]),
      operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1) & and_dcpl_661;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 & and_dcpl_661;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_5_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1,
      nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_4_mux_2_mx0w2,
      nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_5_mux_2_mx0w3,
      {weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_42_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      , and_dcpl_662 , and_dcpl_665});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1,
      operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1, {weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse
      , and_dcpl_661 , and_dcpl_662 , and_dcpl_665});
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse
      = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      = MUX_s_1_2_2(operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1, weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_cse,
      weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      = weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp
      = weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 | (weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1 | (weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1 | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_tmp,
      weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_tmp
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp
      = Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1 | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1 | (weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_6_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_6_sva_1 | (weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 | (weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]));
  assign operator_7_false_1_operator_7_false_1_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 | (weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]));
  assign weight_read_addrs_0_3_0_lpi_1_dfm_4 = MUX_v_4_2_2(4'b0000, pe_manager_base_weight_sva_mx1_3_0,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_4_false_acc_sdt_sva_1 = conv_u2s_4_5(pe_config_num_manager_sva)
      + 5'b11111;
  assign operator_4_false_acc_sdt_sva_1 = nl_operator_4_false_acc_sdt_sva_1[4:0];
  assign while_and_1129_cse_1 = (~ while_if_and_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_if_and_tmp_1 = PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      = ~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl = start_PopNB_mioi_data_rsc_z_mxwt
      & pe_config_is_valid_sva & start_PopNB_mioi_return_rsc_z_mxwt;
  assign PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl = pe_config_is_zero_first_sva
      & pe_manager_zero_active_sva;
  assign PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl = ~(pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign PECore_UpdateFSM_switch_lp_mux1h_14_nl = MUX1HOT_s_1_4_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl,
      PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl, pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1,
      PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl, {PECore_UpdateFSM_switch_lp_and_7_itm_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_2_1 , PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_5_1});
  assign PECore_UpdateFSM_next_state_0_lpi_1_dfm_4 = PECore_UpdateFSM_switch_lp_mux1h_14_nl
      & PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  assign pe_config_UpdateManagerCounter_if_if_unequal_tmp = pe_config_output_counter_sva
      != (operator_8_false_acc_sdt_sva_1[7:0]);
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      = ~(pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]));
  assign input_write_req_valid_lpi_1_dfm_5 = PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      & PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1 = ~(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign or_718_tmp = ((pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2) | and_dcpl_678;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0,
      or_dcpl_296);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4, nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0,
      or_dcpl_296);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5, nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0,
      or_dcpl_296);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0
      = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6, nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0,
      or_dcpl_296);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0,
      or_dcpl_296);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0,
      or_dcpl_296);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0,
      or_dcpl_296);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1 = and_301_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  assign nl_operator_16_false_acc_sdt_sva_1 = conv_u2s_8_9(pe_manager_num_input_sva)
      + 9'b111111111;
  assign operator_16_false_acc_sdt_sva_1 = nl_operator_16_false_acc_sdt_sva_1[8:0];
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1 = ~((state_mux_1_cse!=2'b00)
      | state_0_sva_mx1);
  assign PECore_UpdateFSM_switch_lp_nor_tmp_1 = ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_6 | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1
      | PECore_RunScale_PECore_RunScale_if_and_1_svs_1 | PECore_PushOutput_PECore_PushOutput_if_and_svs_1);
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp
      = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2) | reg_rva_in_reg_rw_sva_2_cse
      | (~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp!=8'b00000000))) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7])));
  assign PECore_DecodeAxiWrite_switch_lp_or_5_cse_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  assign rva_out_reg_data_63_sva_dfm_7 = PECore_PushAxiRsp_mux_13_itm_1 & rva_in_reg_rw_sva_5;
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_1_0_sva_1 = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]!=2'b00));
  assign input_mem_banks_write_if_for_if_and_stg_1_1_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b01);
  assign input_mem_banks_write_if_for_if_and_stg_1_2_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b10);
  assign input_mem_banks_write_if_for_if_and_stg_1_3_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b11);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign nl_PEManager_15U_GetInputAddr_acc_tmp = input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt
      + (pe_manager_base_input_sva[7:0]);
  assign PEManager_15U_GetInputAddr_acc_tmp = nl_PEManager_15U_GetInputAddr_acc_tmp[7:0];
  assign input_write_addrs_lpi_1_dfm_2 = PEManager_15U_GetInputAddr_acc_tmp & ({{7{PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1}},
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1})
      & ({{7{PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1}}, PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1});
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_257_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_255_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_256_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_254_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_255_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_253_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_254_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_252_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_253_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_251_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_252_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_250_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_251_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_249_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_250_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_248_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_249_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_247_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_248_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_246_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_247_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_245_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_246_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_244_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_245_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_243_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_244_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_242_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_243_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_241_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_242_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_240_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_241_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_239_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_240_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_238_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_239_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_237_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_238_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_236_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_237_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_235_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_236_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_234_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_235_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_233_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_234_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_232_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_233_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_231_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_232_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_230_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_231_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_229_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_230_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_228_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_229_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_227_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_228_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_226_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_227_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_225_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_226_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_224_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_225_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_223_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_224_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_222_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_223_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_221_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_222_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_220_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_221_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_219_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_220_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_218_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_219_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_217_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_218_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_216_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_217_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_215_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_216_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_214_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_215_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_213_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_214_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_212_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_213_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_211_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_212_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_210_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_211_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_209_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_210_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_208_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_209_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_207_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_208_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_206_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_207_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_205_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_206_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_204_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_205_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_203_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_204_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_202_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_203_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_201_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_202_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_200_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_201_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_199_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_200_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_198_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_199_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_197_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_198_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_196_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_197_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_195_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_196_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_194_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_195_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_193_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_194_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_192_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_193_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_191_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_192_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_190_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_191_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_189_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_190_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_188_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_189_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_187_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_188_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_186_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_187_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_185_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_186_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_184_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_185_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_183_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_184_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_182_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_183_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_181_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_182_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_180_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_181_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_179_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_180_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_178_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_179_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_177_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_178_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_176_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_177_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_175_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_176_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_174_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_175_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_173_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_174_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_172_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_173_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_171_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_172_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_170_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_171_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_169_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_170_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_168_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_169_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_167_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_168_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_166_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_167_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_165_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_166_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_164_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_165_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_163_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_164_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_162_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_163_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_161_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_162_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_160_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_161_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_159_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_160_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_158_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_159_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_157_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_158_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_156_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_157_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_155_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_156_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_154_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_155_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_153_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_154_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_152_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_153_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_151_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_152_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_150_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_151_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_149_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_150_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_148_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_149_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_147_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_148_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_146_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_147_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_145_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_146_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_144_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_145_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_143_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_144_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_142_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_143_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_141_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_142_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_140_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_141_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_139_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_140_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_138_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_139_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_137_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_138_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_136_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_137_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_135_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_136_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_134_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_135_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_133_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_134_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_132_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_133_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_131_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_132_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_130_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_131_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_129_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_130_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_128_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_129_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_127_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_128_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_126_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_127_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_125_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_126_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_124_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_125_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_123_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_124_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_122_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_123_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_121_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_122_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_120_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_121_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_119_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_120_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_118_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_119_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_117_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_118_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_116_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_117_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_115_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_116_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_114_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_115_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_113_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_114_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_112_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_113_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_111_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_112_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_110_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_111_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_109_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_110_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_108_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_109_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_107_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_108_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_106_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_107_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_105_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_106_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_104_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_105_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_103_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_104_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_102_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_103_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_101_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_102_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_100_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_101_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_99_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_100_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_98_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_99_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_97_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_98_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_96_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_97_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_95_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_96_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_94_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_95_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_93_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_94_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_92_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_93_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_91_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_92_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_90_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_91_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_89_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_90_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_88_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_89_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_87_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_88_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_86_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_87_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_85_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_86_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_84_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_85_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_83_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_84_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_82_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_83_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_81_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_82_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_80_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_81_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_79_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_80_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_78_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_79_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_77_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_78_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_76_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_77_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_75_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_76_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_74_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_75_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_73_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_74_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_72_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_73_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_71_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_72_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_70_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_71_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_69_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_70_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_68_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_69_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_67_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_68_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_66_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_67_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_65_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_66_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_64_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_65_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_63_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_64_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_62_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_63_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_61_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_62_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_60_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_61_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_59_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_60_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_58_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_59_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_57_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_58_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_56_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_57_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_55_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_56_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_54_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_55_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_53_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_54_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_52_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_53_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_51_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_52_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_50_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_51_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_49_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_50_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_48_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_49_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_47_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_48_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_46_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_47_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_45_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_46_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_44_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_45_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_43_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_44_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_42_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_43_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_41_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_42_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_40_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_41_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_39_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_40_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_38_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_39_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_37_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_38_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_36_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_37_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_35_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_36_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_34_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_35_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_33_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_34_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_32_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_33_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_31_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_32_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_30_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_31_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_29_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_30_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_28_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_29_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_27_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_28_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_26_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_27_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_25_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_26_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_24_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_25_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_23_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_24_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_22_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_23_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_21_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_22_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_20_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_21_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_19_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_20_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_18_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_19_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_17_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_18_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_16_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_17_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_15_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_16_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_14_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_15_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_13_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_14_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_12_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_13_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_11_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_12_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_10_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_11_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_9_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_10_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_8_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_9_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_7_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_8_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_6_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_7_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_5_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_6_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_4_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_5_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_3_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_4_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_2_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_3_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_1_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_2_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1 = ~((input_write_addrs_lpi_1_dfm_2[1:0]!=2'b00));
  assign input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b01);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b10);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b11);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2
      | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_4 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0011);
  assign PECore_DecodeAxiRead_switch_lp_nor_13_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_not_185 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 =
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:1]!=15'b000000000000000));
  assign PECore_PushAxiRsp_if_asn_55 = (~ rva_in_reg_rw_sva_10) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_57 = rva_in_reg_rw_sva_10 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_59 = input_read_req_valid_lpi_1_dfm_1_10 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign weight_mem_run_3_for_5_asn_308 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_310 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_312 = (weight_read_addrs_7_lpi_1_dfm_3_2_0[2])
      & nor_690_cse & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_314 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_316 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_318 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_320 = (weight_read_addrs_5_lpi_1_dfm_3_2_0[2])
      & nor_695_cse & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_322 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_324 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_326 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_328 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b100)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_330 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign PECore_PushAxiRsp_if_asn_61 = (~ rva_in_reg_rw_sva_5) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign PECore_PushAxiRsp_if_asn_63 = rva_in_reg_rw_sva_5 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign PECore_PushAxiRsp_if_asn_65 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_166 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_168 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_172 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_174 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign Arbiter_8U_Roundrobin_pick_1_mux_583_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1304_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_583_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_55_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_584_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1303_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_584_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_54_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_585_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1302_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_585_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_53_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_586_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1301_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_586_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_52_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_587_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1300_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_587_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_51_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_588_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_7_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign while_mux_1299_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_588_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_50_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_589_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1297_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_589_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_48_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_590_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1296_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_590_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_47_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_591_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1295_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_591_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_46_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_592_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1294_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_592_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_45_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_593_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1293_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_593_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_44_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_594_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_6_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign while_mux_1292_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_594_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_43_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1291_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_595_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1290_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_595_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_596_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1289_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_596_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_40_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_597_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1288_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_597_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_39_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_598_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1287_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_598_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_38_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_599_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1286_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_599_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_37_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_600_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1285_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_600_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1284_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_607_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1276_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_607_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_608_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1275_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_608_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_609_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1274_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_609_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_610_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1273_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_610_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_611_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1272_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_611_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_612_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1271_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_612_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1270_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_626_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1254_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_626_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_629_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1251_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_629_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_2_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_630_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1250_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_630_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1249_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_dcpl_4 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
      & while_stage_0_11;
  assign and_dcpl_5 = and_dcpl_4 & (~ rva_in_reg_rw_sva_st_1_9);
  assign and_dcpl_6 = and_dcpl_5 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7
      | input_read_req_valid_lpi_1_dfm_1_9 | rva_in_reg_rw_sva_9));
  assign and_dcpl_22 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)
      & while_stage_0_11;
  assign and_dcpl_25 = while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign and_dcpl_27 = while_stage_0_9 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  assign and_dcpl_28 = while_stage_0_9 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign and_dcpl_30 = while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  assign mux_tmp = MUX_s_1_2_2((~ PECore_RunMac_PECore_RunMac_if_and_svs_st_5), rva_in_reg_rw_sva_st_1_5,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_tmp = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_5);
  assign and_dcpl_43 = while_stage_0_6 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign and_dcpl_44 = while_stage_0_6 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_tmp_2 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1 | rva_in_reg_rw_sva_st_1_4;
  assign not_tmp_33 = ~(while_stage_0_4 & PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign and_679_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  assign and_686_cse = weight_mem_read_arbxbar_arbiters_next_7_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign or_38_cse = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_run_3_for_land_4_lpi_1_dfm_1);
  assign or_tmp_60 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign and_dcpl_74 = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
      & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]));
  assign and_dcpl_80 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_81 = and_dcpl_80 & weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  assign and_dcpl_83 = (and_706_cse | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1)
      & and_dcpl_80;
  assign and_dcpl_84 = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      & and_dcpl_80;
  assign and_dcpl_85 = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      & and_dcpl_80;
  assign and_dcpl_86 = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      & and_dcpl_80;
  assign and_dcpl_87 = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      & and_dcpl_80;
  assign and_dcpl_89 = or_708_cse & and_dcpl_80;
  assign and_dcpl_90 = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse
      & and_dcpl_80;
  assign or_dcpl_59 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4);
  assign nor_226_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]));
  assign nor_227_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]));
  assign nor_228_cse = ~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]));
  assign nor_229_cse = ~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]));
  assign nor_233_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]));
  assign nor_231_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]));
  assign and_107_cse = (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]) |
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]))) & nor_231_cse & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]))) & nor_233_cse;
  assign nor_237_cse = ~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]));
  assign and_114_cse = (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]) |
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]))) & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]))) & nor_237_cse;
  assign and_121_cse = (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]) |
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]))) & (~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])));
  assign nor_242_cse = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]));
  assign and_128_cse = nor_242_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])));
  assign nor_246_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]));
  assign and_135_cse = nor_246_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])));
  assign nor_253_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]));
  assign and_142_cse = (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) |
      (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]))) & nor_253_cse;
  assign or_dcpl_68 = and_142_cse | or_dcpl_59;
  assign and_dcpl_140 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign and_dcpl_141 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign and_dcpl_142 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign and_dcpl_143 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign and_dcpl_144 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign and_dcpl_145 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign and_dcpl_146 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign and_dcpl_147 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign and_dcpl_153 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_158 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign and_dcpl_170 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_171 = and_dcpl_144 & and_dcpl_153;
  assign and_dcpl_173 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_174 = and_dcpl_143 & and_dcpl_153;
  assign and_dcpl_176 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_177 = and_dcpl_145 & and_dcpl_153;
  assign and_dcpl_179 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_180 = and_dcpl_147 & and_dcpl_153;
  assign and_dcpl_182 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_183 = and_dcpl_141 & and_dcpl_153;
  assign and_dcpl_185 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_186 = and_dcpl_142 & and_dcpl_153;
  assign and_dcpl_187 = and_dcpl_153 & (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]);
  assign and_dcpl_188 = and_dcpl_153 & and_dcpl_140;
  assign and_dcpl_190 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_191 = and_dcpl_146 & and_dcpl_153;
  assign and_dcpl_194 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign and_dcpl_198 = (state_2_1_sva==2'b01) & (~ state_0_sva) & and_604_cse;
  assign mux_41_nl = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      state_2_1_sva[1]);
  assign and_699_nl = (state_2_1_sva[1]) & PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  assign mux_42_nl = MUX_s_1_2_2(mux_41_nl, and_699_nl, state_2_1_sva[0]);
  assign mux_43_nl = MUX_s_1_2_2(mux_42_nl, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      state_0_sva);
  assign and_dcpl_201 = mux_43_nl & (~(PECore_RunFSM_switch_lp_nor_tmp_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign or_dcpl_135 = ~(rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse);
  assign or_dcpl_141 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]!=2'b01);
  assign and_dcpl_203 = reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign and_dcpl_206 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01);
  assign and_dcpl_207 = and_dcpl_206 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]))
      & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign and_dcpl_208 = and_dcpl_207 & and_dcpl_203 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_209 = reg_rva_in_PopNB_mioi_iswt0_cse & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_211 = and_dcpl_207 & and_dcpl_209 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign or_tmp_84 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1 |
      rva_in_reg_rw_sva_st_1_4 | rva_in_reg_rw_sva_4;
  assign mux_59_nl = MUX_s_1_2_2((~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])),
      (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_tmp_60 = MUX_s_1_2_2(mux_59_nl, or_231_cse, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign or_238_nl = (~((~((~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign or_234_nl = (~((~((~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign mux_tmp_62 = MUX_s_1_2_2(or_238_nl, or_234_nl, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_tmp_94 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | mux_tmp_62;
  assign or_tmp_95 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ mux_tmp_62);
  assign nor_260_cse = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2:1]!=2'b00));
  assign and_dcpl_240 = rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign and_dcpl_244 = while_stage_0_10 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  assign and_dcpl_245 = and_dcpl_240 & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_248 = PECore_RunFSM_switch_lp_equal_tmp_1_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_267 = and_dcpl_244 & (~ rva_in_reg_rw_sva_st_1_8);
  assign or_tmp_111 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_run_3_for_weight_mem_run_3_for_and_4_cse);
  assign and_dcpl_284 = and_dcpl_267 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6
      | rva_in_reg_rw_sva_8 | input_read_req_valid_lpi_1_dfm_1_8));
  assign and_dcpl_297 = and_dcpl_206 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]))
      & and_dcpl_240;
  assign and_dcpl_305 = and_dcpl_27 & (~ rva_in_reg_rw_sva_st_1_7);
  assign and_dcpl_308 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5
      | rva_in_reg_rw_sva_7 | input_read_req_valid_lpi_1_dfm_1_7);
  assign and_dcpl_309 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & (~ rva_in_reg_rw_sva_st_1_7);
  assign not_tmp_182 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1
      | reg_rva_in_reg_rw_sva_2_cse);
  assign and_dcpl_325 = and_dcpl_30 & (~ rva_in_reg_rw_sva_st_1_6);
  assign and_dcpl_337 = and_dcpl_325 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4
      | rva_in_reg_rw_sva_6 | input_read_req_valid_lpi_1_dfm_1_6));
  assign and_dcpl_349 = (~ rva_in_reg_rw_sva_st_1_5) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign and_dcpl_350 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | rva_in_reg_rw_sva_5);
  assign and_dcpl_357 = and_dcpl_349 & while_stage_0_7;
  assign and_dcpl_375 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7;
  assign and_dcpl_393 = ~(rva_in_reg_rw_sva_st_1_3 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1);
  assign and_dcpl_406 = and_dcpl_393 & (~ input_read_req_valid_lpi_1_dfm_1_3);
  assign and_dcpl_417 = (crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_1_tmp | (~
      weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp))
      & (~(reg_rva_in_reg_rw_sva_2_cse | input_read_req_valid_lpi_1_dfm_1_2));
  assign and_dcpl_434 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | input_read_req_valid_lpi_1_dfm_1_1);
  assign and_dcpl_435 = and_dcpl_434 & and_dcpl_194;
  assign mux_tmp_97 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1!=4'b0100));
  assign and_dcpl_441 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1);
  assign nand_31_cse = ~(PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]));
  assign and_dcpl_476 = PECore_RunMac_PECore_RunMac_if_and_svs_st_7 & while_stage_0_9
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign and_dcpl_480 = while_stage_0_8 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
  assign and_dcpl_486 = (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign mux_tmp_98 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_496_nl = while_stage_0_6 & mux_tmp_98;
  assign and_495_nl = while_stage_0_6 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_tmp_99 = MUX_s_1_2_2(and_496_nl, and_495_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1);
  assign and_dcpl_489 = and_882_cse & (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign mux_tmp_102 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_501_nl = while_stage_0_6 & mux_tmp_102;
  assign and_500_nl = while_stage_0_6 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_tmp_103 = MUX_s_1_2_2(and_501_nl, and_500_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1);
  assign nor_320_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1);
  assign mux_106_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_320_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign not_tmp_264 = while_stage_0_6 & mux_106_nl;
  assign nor_321_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1);
  assign mux_108_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_321_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign not_tmp_267 = while_stage_0_6 & mux_108_nl;
  assign and_719_nl = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & while_stage_0_6;
  assign nor_322_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1 | (~ while_stage_0_6));
  assign not_tmp_270 = MUX_s_1_2_2(and_719_nl, nor_322_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_tmp_164 = (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1 | (~ while_stage_0_6);
  assign nor_tmp_47 = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & while_stage_0_6;
  assign or_374_nl = while_stage_0_5 | nor_tmp_47;
  assign or_373_nl = while_stage_0_5 | (~ or_tmp_164);
  assign mux_tmp_113 = MUX_s_1_2_2(or_374_nl, or_373_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign not_tmp_274 = MUX_s_1_2_2(nor_tmp_47, (~ or_tmp_164), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_722_nl = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & while_stage_0_6;
  assign nor_323_nl = ~((~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1 | (~ while_stage_0_6));
  assign not_tmp_277 = MUX_s_1_2_2(and_722_nl, nor_323_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_tmp_178 = (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1 | (~ while_stage_0_6);
  assign nor_tmp_50 = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & while_stage_0_6;
  assign or_390_nl = while_stage_0_5 | nor_tmp_50;
  assign or_389_nl = while_stage_0_5 | (~ or_tmp_178);
  assign mux_tmp_123 = MUX_s_1_2_2(or_390_nl, or_389_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign not_tmp_281 = MUX_s_1_2_2(nor_tmp_50, (~ or_tmp_178), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_dcpl_218 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7);
  assign and_dcpl_543 = nor_226_cse & nor_227_cse;
  assign and_dcpl_544 = and_dcpl_543 & nor_228_cse & nor_229_cse;
  assign and_dcpl_545 = and_dcpl_80 & (~ while_stage_0_4);
  assign or_dcpl_227 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ while_stage_0_5);
  assign or_dcpl_228 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ while_stage_0_3);
  assign or_dcpl_239 = or_dcpl_135 | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_240 = or_dcpl_141 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]);
  assign and_dcpl_594 = nor_260_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign and_dcpl_595 = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign and_dcpl_596 = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2:1]==2'b10);
  assign and_dcpl_597 = and_dcpl_596 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign and_dcpl_599 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]));
  assign and_dcpl_603 = ~(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_dcpl_275 = (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | nand_31_cse;
  assign or_dcpl_278 = PECore_RunMac_PECore_RunMac_if_and_svs_st_8 | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_8);
  assign or_dcpl_283 = (~(while_stage_0_8 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6))
      | rva_in_reg_rw_sva_6;
  assign nor_tmp_58 = while_mux_1299_tmp & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign and_728_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) & while_mux_1300_tmp;
  assign while_mux_1298_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_206 = and_728_cse | while_mux_1298_nl | nor_tmp_58;
  assign or_495_nl = and_728_cse | nor_tmp_58;
  assign mux_tmp_152 = MUX_s_1_2_2(or_495_nl, or_tmp_206, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign or_tmp_208 = and_679_cse | and_686_cse;
  assign or_tmp_209 = ((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1)
      | or_tmp_208;
  assign mux_tmp_153 = MUX_s_1_2_2(or_tmp_209, mux_tmp_152, while_stage_0_5);
  assign nand_8_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      & (~ or_tmp_209));
  assign mux_157_nl = MUX_s_1_2_2(nand_8_nl, or_tmp_209, and_889_cse);
  assign mux_158_nl = MUX_s_1_2_2(mux_157_nl, or_tmp_209, and_888_cse);
  assign mux_159_nl = MUX_s_1_2_2(mux_158_nl, or_tmp_209, and_887_cse);
  assign nand_7_nl = ~(while_mux_1302_tmp & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      & (~ mux_tmp_152));
  assign mux_154_nl = MUX_s_1_2_2(nand_7_nl, mux_tmp_152, and_893_cse);
  assign mux_155_nl = MUX_s_1_2_2(mux_154_nl, mux_tmp_152, and_892_cse);
  assign mux_156_nl = MUX_s_1_2_2(mux_155_nl, mux_tmp_152, and_891_cse);
  assign mux_160_itm = MUX_s_1_2_2(mux_159_nl, mux_156_nl, while_stage_0_5);
  assign or_506_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]));
  assign mux_164_nl = MUX_s_1_2_2(or_506_nl, and_686_cse, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign or_505_nl = weight_mem_read_arbxbar_arbiters_next_7_5_sva | and_686_cse;
  assign mux_165_nl = MUX_s_1_2_2(mux_164_nl, or_505_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign or_504_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | or_tmp_208;
  assign mux_166_nl = MUX_s_1_2_2(mux_165_nl, or_504_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign nor_358_nl = ~(and_887_cse | and_888_cse | and_889_cse | and_890_cse | mux_166_nl);
  assign or_499_nl = while_mux_1299_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]));
  assign mux_161_nl = MUX_s_1_2_2(or_499_nl, nor_tmp_58, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign or_498_nl = while_mux_1300_tmp | nor_tmp_58;
  assign mux_162_nl = MUX_s_1_2_2(mux_161_nl, or_498_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign mux_163_nl = MUX_s_1_2_2(mux_162_nl, or_tmp_206, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign nor_359_nl = ~(and_891_cse | and_892_cse | and_893_cse | and_894_cse | mux_163_nl);
  assign not_tmp_425 = MUX_s_1_2_2(nor_358_nl, nor_359_nl, while_stage_0_5);
  assign or_tmp_223 = and_893_cse | and_894_cse;
  assign or_tmp_229 = and_889_cse | and_890_cse;
  assign nor_360_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_3_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])));
  assign nor_361_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_2_sva | and_890_cse);
  assign mux_171_nl = MUX_s_1_2_2(nor_360_nl, nor_361_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign nor_362_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_4_sva | or_tmp_229);
  assign mux_172_nl = MUX_s_1_2_2(mux_171_nl, nor_362_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign nor_363_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_1_sva | and_888_cse
      | or_tmp_229);
  assign mux_173_nl = MUX_s_1_2_2(mux_172_nl, nor_363_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign nor_364_nl = ~(while_mux_1302_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])));
  assign nor_365_nl = ~(while_mux_1303_tmp | and_894_cse);
  assign mux_168_nl = MUX_s_1_2_2(nor_364_nl, nor_365_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign nor_366_nl = ~(while_mux_1301_tmp | or_tmp_223);
  assign mux_169_nl = MUX_s_1_2_2(mux_168_nl, nor_366_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign nor_367_nl = ~(while_mux_1304_tmp | and_892_cse | or_tmp_223);
  assign mux_170_nl = MUX_s_1_2_2(mux_169_nl, nor_367_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign mux_174_nl = MUX_s_1_2_2(mux_173_nl, mux_170_nl, while_stage_0_5);
  assign and_dcpl_632 = mux_174_nl & and_dcpl_543;
  assign and_755_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & while_mux_1293_tmp;
  assign and_756_cse = while_mux_1292_tmp & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign or_tmp_243 = and_755_cse | and_756_cse;
  assign and_757_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  assign and_758_cse = weight_mem_read_arbxbar_arbiters_next_6_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign or_tmp_245 = and_757_cse | and_758_cse;
  assign mux_177_nl = MUX_s_1_2_2(or_tmp_245, or_tmp_243, while_stage_0_5);
  assign or_534_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | or_tmp_245;
  assign or_532_nl = while_mux_1291_tmp | or_tmp_243;
  assign mux_176_nl = MUX_s_1_2_2(or_534_nl, or_532_nl, while_stage_0_5);
  assign mux_tmp_178 = MUX_s_1_2_2(mux_177_nl, mux_176_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_tmp_247 = while_mux_1295_tmp | while_mux_1297_tmp;
  assign and_761_cse = while_mux_1291_tmp & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_tmp_249 = and_755_cse | and_756_cse | and_761_cse;
  assign and_763_cse = while_mux_1296_tmp & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign or_tmp_250 = weight_mem_read_arbxbar_arbiters_next_6_3_sva | weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  assign or_tmp_252 = and_757_cse | and_758_cse | ((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1);
  assign and_768_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  assign nand_10_nl = ~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_4_sva
      & (~ or_tmp_252));
  assign mux_181_itm = MUX_s_1_2_2(nand_10_nl, or_tmp_252, and_768_cse);
  assign nand_9_nl = ~(while_mux_1294_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      & (~ or_tmp_249));
  assign mux_179_itm = MUX_s_1_2_2(nand_9_nl, or_tmp_249, and_763_cse);
  assign mux_191_nl = MUX_s_1_2_2(mux_181_itm, mux_179_itm, while_stage_0_5);
  assign mux_189_nl = MUX_s_1_2_2(mux_181_itm, or_tmp_252, weight_mem_read_arbxbar_arbiters_next_6_3_sva);
  assign mux_188_nl = MUX_s_1_2_2(mux_179_itm, or_tmp_249, while_mux_1295_tmp);
  assign mux_190_nl = MUX_s_1_2_2(mux_189_nl, mux_188_nl, while_stage_0_5);
  assign mux_192_nl = MUX_s_1_2_2(mux_191_nl, mux_190_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_185_nl = MUX_s_1_2_2(mux_181_itm, or_tmp_252, weight_mem_read_arbxbar_arbiters_next_6_1_sva);
  assign mux_184_nl = MUX_s_1_2_2(mux_179_itm, or_tmp_249, while_mux_1297_tmp);
  assign mux_186_nl = MUX_s_1_2_2(mux_185_nl, mux_184_nl, while_stage_0_5);
  assign mux_182_nl = MUX_s_1_2_2(mux_181_itm, or_tmp_252, or_tmp_250);
  assign mux_180_nl = MUX_s_1_2_2(mux_179_itm, or_tmp_249, or_tmp_247);
  assign mux_183_nl = MUX_s_1_2_2(mux_182_nl, mux_180_nl, while_stage_0_5);
  assign mux_187_nl = MUX_s_1_2_2(mux_186_nl, mux_183_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_193_itm = MUX_s_1_2_2(mux_192_nl, mux_187_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_tmp_254 = and_761_cse | and_756_cse;
  assign and_772_cse = while_mux_1294_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign or_545_nl = while_mux_1292_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign or_544_nl = while_mux_1291_tmp | and_756_cse;
  assign mux_194_nl = MUX_s_1_2_2(or_545_nl, or_544_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_195_nl = MUX_s_1_2_2(mux_194_nl, or_tmp_254, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_543_nl = while_mux_1293_tmp | or_tmp_254;
  assign mux_196_nl = MUX_s_1_2_2(mux_195_nl, or_543_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_259 = and_763_cse | and_772_cse | mux_196_nl;
  assign or_tmp_262 = and_758_cse | Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  assign mux_tmp_197 = MUX_s_1_2_2(and_758_cse, or_tmp_262, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign and_776_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  assign or_552_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign mux_198_nl = MUX_s_1_2_2(or_552_nl, or_tmp_262, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign mux_199_nl = MUX_s_1_2_2(mux_198_nl, mux_tmp_197, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign or_551_nl = weight_mem_read_arbxbar_arbiters_next_6_5_sva | mux_tmp_197;
  assign mux_200_nl = MUX_s_1_2_2(mux_199_nl, or_551_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign or_tmp_266 = and_768_cse | and_776_cse | mux_200_nl;
  assign mux_205_nl = MUX_s_1_2_2(or_tmp_266, or_tmp_259, while_stage_0_5);
  assign or_559_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | or_tmp_266;
  assign or_558_nl = while_mux_1295_tmp | or_tmp_259;
  assign mux_204_nl = MUX_s_1_2_2(or_559_nl, or_558_nl, while_stage_0_5);
  assign mux_206_nl = MUX_s_1_2_2(mux_205_nl, mux_204_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign or_557_nl = weight_mem_read_arbxbar_arbiters_next_6_1_sva | or_tmp_266;
  assign or_556_nl = while_mux_1297_tmp | or_tmp_259;
  assign mux_202_nl = MUX_s_1_2_2(or_557_nl, or_556_nl, while_stage_0_5);
  assign or_555_nl = or_tmp_250 | or_tmp_266;
  assign or_548_nl = or_tmp_247 | or_tmp_259;
  assign mux_201_nl = MUX_s_1_2_2(or_555_nl, or_548_nl, while_stage_0_5);
  assign mux_203_nl = MUX_s_1_2_2(mux_202_nl, mux_201_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_207_itm = MUX_s_1_2_2(mux_206_nl, mux_203_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign nor_tmp_117 = while_mux_1297_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_tmp_272 = and_763_cse | nor_tmp_117;
  assign nor_tmp_120 = weight_mem_read_arbxbar_arbiters_next_6_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_tmp_278 = and_768_cse | nor_tmp_120;
  assign and_782_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & while_mux_1295_tmp;
  assign and_781_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  assign nor_368_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_1_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])));
  assign nor_369_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_2_sva | nor_tmp_120);
  assign mux_211_nl = MUX_s_1_2_2(nor_368_nl, nor_369_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign nor_370_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_3_sva | or_tmp_278);
  assign mux_212_nl = MUX_s_1_2_2(mux_211_nl, nor_370_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nor_371_nl = ~(weight_mem_read_arbxbar_arbiters_next_6_4_sva | and_781_cse
      | or_tmp_278);
  assign mux_213_nl = MUX_s_1_2_2(mux_212_nl, nor_371_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign nor_372_nl = ~(while_mux_1297_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])));
  assign nor_373_nl = ~(while_mux_1296_tmp | nor_tmp_117);
  assign mux_208_nl = MUX_s_1_2_2(nor_372_nl, nor_373_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign nor_374_nl = ~(while_mux_1295_tmp | or_tmp_272);
  assign mux_209_nl = MUX_s_1_2_2(mux_208_nl, nor_374_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nor_375_nl = ~(while_mux_1294_tmp | and_782_cse | or_tmp_272);
  assign mux_210_nl = MUX_s_1_2_2(mux_209_nl, nor_375_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign mux_214_nl = MUX_s_1_2_2(mux_213_nl, mux_210_nl, while_stage_0_5);
  assign and_dcpl_634 = mux_214_nl & nor_231_cse & nor_233_cse;
  assign or_tmp_287 = and_772_cse | and_782_cse | and_755_cse | and_756_cse | or_tmp_272;
  assign or_tmp_292 = and_776_cse | and_781_cse | and_757_cse | and_758_cse | or_tmp_278;
  assign and_792_cse = while_mux_1286_tmp & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign and_791_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) & while_mux_1285_tmp;
  assign or_tmp_294 = and_791_cse | and_792_cse;
  assign and_794_cse = weight_mem_read_arbxbar_arbiters_next_5_5_sva & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign and_793_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  assign or_tmp_296 = and_793_cse | and_794_cse;
  assign mux_219_nl = MUX_s_1_2_2(or_tmp_296, or_tmp_294, while_stage_0_5);
  assign or_585_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1
      | or_tmp_296;
  assign or_583_nl = while_mux_1284_tmp | or_tmp_294;
  assign mux_218_nl = MUX_s_1_2_2(or_585_nl, or_583_nl, while_stage_0_5);
  assign mux_tmp_220 = MUX_s_1_2_2(mux_219_nl, mux_218_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign or_tmp_300 = and_792_cse | and_791_cse | (while_mux_1284_tmp & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]));
  assign or_tmp_303 = and_794_cse | and_793_cse | ((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1);
  assign and_804_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  assign nand_12_nl = ~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_4_sva
      & (~ or_tmp_303));
  assign mux_223_itm = MUX_s_1_2_2(nand_12_nl, or_tmp_303, and_804_cse);
  assign nand_11_nl = ~(while_mux_1287_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      & (~ or_tmp_300));
  assign and_799_nl = while_mux_1289_tmp & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign mux_221_itm = MUX_s_1_2_2(nand_11_nl, or_tmp_300, and_799_nl);
  assign mux_233_nl = MUX_s_1_2_2(mux_223_itm, mux_221_itm, while_stage_0_5);
  assign mux_231_nl = MUX_s_1_2_2(mux_223_itm, or_tmp_303, weight_mem_read_arbxbar_arbiters_next_5_3_sva);
  assign mux_230_nl = MUX_s_1_2_2(mux_221_itm, or_tmp_300, while_mux_1288_tmp);
  assign mux_232_nl = MUX_s_1_2_2(mux_231_nl, mux_230_nl, while_stage_0_5);
  assign mux_234_nl = MUX_s_1_2_2(mux_233_nl, mux_232_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign mux_227_nl = MUX_s_1_2_2(mux_223_itm, or_tmp_303, weight_mem_read_arbxbar_arbiters_next_5_1_sva);
  assign mux_226_nl = MUX_s_1_2_2(mux_221_itm, or_tmp_300, while_mux_1290_tmp);
  assign mux_228_nl = MUX_s_1_2_2(mux_227_nl, mux_226_nl, while_stage_0_5);
  assign or_589_nl = weight_mem_read_arbxbar_arbiters_next_5_3_sva | weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  assign mux_224_nl = MUX_s_1_2_2(mux_223_itm, or_tmp_303, or_589_nl);
  assign or_586_nl = while_mux_1288_tmp | while_mux_1290_tmp;
  assign mux_222_nl = MUX_s_1_2_2(mux_221_itm, or_tmp_300, or_586_nl);
  assign mux_225_nl = MUX_s_1_2_2(mux_224_nl, mux_222_nl, while_stage_0_5);
  assign mux_229_nl = MUX_s_1_2_2(mux_228_nl, mux_225_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign mux_235_itm = MUX_s_1_2_2(mux_234_nl, mux_229_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign and_805_cse = while_mux_1290_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign or_tmp_304 = and_805_cse | while_mux_1289_tmp;
  assign mux_tmp_236 = MUX_s_1_2_2(and_805_cse, or_tmp_304, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign or_tmp_305 = ((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]) & while_mux_1288_tmp)
      | mux_tmp_236;
  assign or_tmp_306 = and_792_cse | or_tmp_305;
  assign and_809_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) & while_mux_1287_tmp;
  assign or_tmp_308 = and_809_cse | and_791_cse | or_tmp_306;
  assign nor_tmp_154 = weight_mem_read_arbxbar_arbiters_next_5_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]);
  assign or_tmp_310 = and_804_cse | nor_tmp_154;
  assign or_tmp_311 = ((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_3_sva)
      | or_tmp_310;
  assign or_tmp_312 = and_794_cse | or_tmp_311;
  assign and_815_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  assign or_tmp_314 = and_815_cse | and_793_cse | or_tmp_312;
  assign or_603_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1
      | or_tmp_314;
  assign or_597_nl = while_mux_1284_tmp | or_tmp_308;
  assign mux_tmp_237 = MUX_s_1_2_2(or_603_nl, or_597_nl, while_stage_0_5);
  assign mux_238_nl = MUX_s_1_2_2(or_tmp_314, or_tmp_308, while_stage_0_5);
  assign mux_tmp_239 = MUX_s_1_2_2(mux_238_nl, mux_tmp_237, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign or_701_nl = weight_mem_read_arbxbar_arbiters_next_5_5_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]))
      | or_tmp_311;
  assign or_606_nl = weight_mem_read_arbxbar_arbiters_next_5_6_sva | or_tmp_312;
  assign mux_241_nl = MUX_s_1_2_2(or_701_nl, or_606_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign or_607_nl = and_815_cse | mux_241_nl;
  assign or_702_nl = while_mux_1286_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]))
      | or_tmp_305;
  assign or_604_nl = while_mux_1285_tmp | or_tmp_306;
  assign mux_240_nl = MUX_s_1_2_2(or_702_nl, or_604_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign or_605_nl = and_809_cse | mux_240_nl;
  assign mux_242_nl = MUX_s_1_2_2(or_607_nl, or_605_nl, while_stage_0_5);
  assign mux_243_nl = MUX_s_1_2_2(mux_242_nl, mux_tmp_237, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign mux_244_itm = MUX_s_1_2_2(mux_243_nl, mux_tmp_239, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign or_614_nl = weight_mem_read_arbxbar_arbiters_next_5_1_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]));
  assign or_613_nl = weight_mem_read_arbxbar_arbiters_next_5_2_sva | nor_tmp_154;
  assign mux_248_nl = MUX_s_1_2_2(or_614_nl, or_613_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign or_612_nl = weight_mem_read_arbxbar_arbiters_next_5_3_sva | or_tmp_310;
  assign mux_249_nl = MUX_s_1_2_2(mux_248_nl, or_612_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign or_611_nl = weight_mem_read_arbxbar_arbiters_next_5_4_sva | or_tmp_311;
  assign mux_250_nl = MUX_s_1_2_2(mux_249_nl, or_611_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign or_610_nl = while_mux_1290_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]));
  assign mux_245_nl = MUX_s_1_2_2(or_610_nl, or_tmp_304, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign or_609_nl = while_mux_1288_tmp | mux_tmp_236;
  assign mux_246_nl = MUX_s_1_2_2(mux_245_nl, or_609_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign or_608_nl = while_mux_1287_tmp | or_tmp_305;
  assign mux_247_nl = MUX_s_1_2_2(mux_246_nl, or_608_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign mux_251_nl = MUX_s_1_2_2(mux_250_nl, mux_247_nl, while_stage_0_5);
  assign and_dcpl_637 = (~ mux_251_nl) & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]))) & nor_237_cse;
  assign while_mux_1277_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_252 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1,
      while_mux_1277_nl, while_stage_0_5);
  assign and_dcpl_639 = (mux_tmp_252 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]))
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp;
  assign and_dcpl_642 = (~(mux_tmp_252 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])))
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp))
      & weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp;
  assign and_dcpl_643 = weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_dcpl_644 = ~(weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_5_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_820_cse = while_mux_1271_tmp & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign or_tmp_327 = ((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]) & while_mux_1272_tmp)
      | and_820_cse;
  assign and_822_cse = weight_mem_read_arbxbar_arbiters_next_3_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign or_tmp_329 = ((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_5_sva)
      | and_822_cse;
  assign mux_254_nl = MUX_s_1_2_2(or_tmp_329, or_tmp_327, while_stage_0_5);
  assign or_621_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1
      | or_tmp_329;
  assign or_619_nl = while_mux_1270_tmp | or_tmp_327;
  assign mux_253_nl = MUX_s_1_2_2(or_621_nl, or_619_nl, while_stage_0_5);
  assign mux_tmp_255 = MUX_s_1_2_2(mux_254_nl, mux_253_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign and_824_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) & while_mux_1275_tmp;
  assign and_825_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) & while_mux_1273_tmp;
  assign and_826_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]) & while_mux_1274_tmp;
  assign nand_15_nl = ~(while_mux_1276_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])
      & (~ or_tmp_327));
  assign mux_256_nl = MUX_s_1_2_2(nand_15_nl, or_tmp_327, and_824_cse);
  assign mux_257_nl = MUX_s_1_2_2(mux_256_nl, or_tmp_327, and_825_cse);
  assign mux_tmp_258 = MUX_s_1_2_2(mux_257_nl, or_tmp_327, and_826_cse);
  assign and_828_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  assign and_829_cse = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_4_sva;
  assign and_830_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  assign nand_16_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])
      & (~ or_tmp_329));
  assign mux_259_nl = MUX_s_1_2_2(nand_16_nl, or_tmp_329, and_828_cse);
  assign mux_260_nl = MUX_s_1_2_2(mux_259_nl, or_tmp_329, and_829_cse);
  assign mux_tmp_261 = MUX_s_1_2_2(mux_260_nl, or_tmp_329, and_830_cse);
  assign mux_263_nl = MUX_s_1_2_2(mux_tmp_261, mux_tmp_258, while_stage_0_5);
  assign or_623_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1
      | mux_tmp_261;
  assign or_622_nl = while_mux_1270_tmp | mux_tmp_258;
  assign mux_262_nl = MUX_s_1_2_2(or_623_nl, or_622_nl, while_stage_0_5);
  assign mux_264_itm = MUX_s_1_2_2(mux_263_nl, mux_262_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign or_tmp_334 = ((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]) & while_mux_1270_tmp)
      | and_820_cse;
  assign or_628_nl = while_mux_1271_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]));
  assign or_627_nl = while_mux_1270_tmp | and_820_cse;
  assign mux_265_nl = MUX_s_1_2_2(or_628_nl, or_627_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign mux_266_nl = MUX_s_1_2_2(mux_265_nl, or_tmp_334, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign or_626_nl = while_mux_1272_tmp | or_tmp_334;
  assign mux_267_nl = MUX_s_1_2_2(mux_266_nl, or_626_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign or_tmp_339 = and_824_cse | and_825_cse | mux_267_nl;
  assign or_tmp_342 = ((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1)
      | and_822_cse;
  assign or_636_nl = weight_mem_read_arbxbar_arbiters_next_3_6_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]));
  assign or_635_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1
      | and_822_cse;
  assign mux_268_nl = MUX_s_1_2_2(or_636_nl, or_635_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign mux_269_nl = MUX_s_1_2_2(mux_268_nl, or_tmp_342, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign or_634_nl = weight_mem_read_arbxbar_arbiters_next_3_5_sva | or_tmp_342;
  assign mux_270_nl = MUX_s_1_2_2(mux_269_nl, or_634_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign or_tmp_347 = and_828_cse | and_829_cse | mux_270_nl;
  assign mux_275_nl = MUX_s_1_2_2(or_tmp_347, or_tmp_339, while_stage_0_5);
  assign or_643_nl = weight_mem_read_arbxbar_arbiters_next_3_3_sva | or_tmp_347;
  assign or_642_nl = while_mux_1274_tmp | or_tmp_339;
  assign mux_274_nl = MUX_s_1_2_2(or_643_nl, or_642_nl, while_stage_0_5);
  assign mux_276_nl = MUX_s_1_2_2(mux_275_nl, mux_274_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign or_641_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva | or_tmp_347;
  assign or_640_nl = while_mux_1276_tmp | or_tmp_339;
  assign mux_272_nl = MUX_s_1_2_2(or_641_nl, or_640_nl, while_stage_0_5);
  assign or_639_nl = weight_mem_read_arbxbar_arbiters_next_3_1_sva | weight_mem_read_arbxbar_arbiters_next_3_3_sva
      | or_tmp_347;
  assign or_631_nl = while_mux_1274_tmp | while_mux_1276_tmp | or_tmp_339;
  assign mux_271_nl = MUX_s_1_2_2(or_639_nl, or_631_nl, while_stage_0_5);
  assign mux_273_nl = MUX_s_1_2_2(mux_272_nl, mux_271_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign mux_277_itm = MUX_s_1_2_2(mux_276_nl, mux_273_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign nor_tmp_181 = while_mux_1276_tmp & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign or_tmp_353 = and_824_cse | nor_tmp_181;
  assign nor_tmp_184 = weight_mem_read_arbxbar_arbiters_next_3_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign or_tmp_359 = and_828_cse | nor_tmp_184;
  assign nor_379_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_1_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])));
  assign nor_380_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_2_sva | nor_tmp_184);
  assign mux_281_nl = MUX_s_1_2_2(nor_379_nl, nor_380_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign nor_381_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_4_sva | or_tmp_359);
  assign mux_282_nl = MUX_s_1_2_2(mux_281_nl, nor_381_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign nor_382_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_3_sva | and_829_cse
      | or_tmp_359);
  assign mux_283_nl = MUX_s_1_2_2(mux_282_nl, nor_382_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign nor_383_nl = ~(while_mux_1276_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])));
  assign nor_384_nl = ~(while_mux_1275_tmp | nor_tmp_181);
  assign mux_278_nl = MUX_s_1_2_2(nor_383_nl, nor_384_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign nor_385_nl = ~(while_mux_1273_tmp | or_tmp_353);
  assign mux_279_nl = MUX_s_1_2_2(mux_278_nl, nor_385_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign nor_386_nl = ~(while_mux_1274_tmp | and_825_cse | or_tmp_353);
  assign mux_280_nl = MUX_s_1_2_2(mux_279_nl, nor_386_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign mux_284_nl = MUX_s_1_2_2(mux_283_nl, mux_280_nl, while_stage_0_5);
  assign and_dcpl_647 = mux_284_nl & nor_242_cse & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])));
  assign or_tmp_368 = and_826_cse | and_825_cse | and_824_cse | nor_tmp_181 | or_tmp_327;
  assign or_tmp_373 = and_830_cse | and_829_cse | and_828_cse | nor_tmp_184 | or_tmp_329;
  assign and_853_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) & while_mux_1250_tmp;
  assign and_854_cse = while_mux_1251_tmp & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign or_tmp_375 = and_853_cse | and_854_cse;
  assign and_855_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) & weight_mem_read_arbxbar_arbiters_next_0_6_sva;
  assign and_856_cse = weight_mem_read_arbxbar_arbiters_next_0_5_sva & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign or_tmp_377 = and_855_cse | and_856_cse;
  assign mux_289_nl = MUX_s_1_2_2(or_tmp_377, or_tmp_375, while_stage_0_5);
  assign or_669_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | or_tmp_377;
  assign or_667_nl = while_mux_1249_tmp | or_tmp_375;
  assign mux_288_nl = MUX_s_1_2_2(or_669_nl, or_667_nl, while_stage_0_5);
  assign mux_tmp_290 = MUX_s_1_2_2(mux_289_nl, mux_288_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign or_tmp_379 = weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_mux_625_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1255_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_625_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_859_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]) & while_mux_1255_nl;
  assign Arbiter_8U_Roundrobin_pick_1_mux_627_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1253_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_627_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_4_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_860_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]) & while_mux_1253_nl;
  assign mux_291_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp,
      or_tmp_379, while_mux_1254_tmp);
  assign or_tmp_383 = and_853_cse | and_854_cse | (~(and_859_cse | and_860_cse |
      mux_291_nl));
  assign and_863_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]) & weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  assign and_864_cse = weight_mem_read_arbxbar_arbiters_next_0_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign mux_292_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp,
      or_tmp_379, weight_mem_read_arbxbar_arbiters_next_0_2_sva);
  assign or_tmp_388 = and_855_cse | and_856_cse | (~(and_863_cse | and_864_cse |
      mux_292_nl));
  assign mux_294_nl = MUX_s_1_2_2(or_tmp_388, or_tmp_383, while_stage_0_5);
  assign or_680_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | or_tmp_388;
  assign or_675_nl = while_mux_1249_tmp | or_tmp_383;
  assign mux_293_nl = MUX_s_1_2_2(or_680_nl, or_675_nl, while_stage_0_5);
  assign mux_295_itm = MUX_s_1_2_2(mux_294_nl, mux_293_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign or_tmp_391 = and_859_cse | and_860_cse | (while_mux_1254_tmp & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]));
  assign or_tmp_392 = and_854_cse | or_tmp_391;
  assign or_tmp_393 = and_853_cse | or_tmp_392;
  assign or_tmp_396 = and_863_cse | and_864_cse | (weight_mem_read_arbxbar_arbiters_next_0_2_sva
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]));
  assign or_tmp_397 = and_856_cse | or_tmp_396;
  assign or_tmp_398 = and_855_cse | or_tmp_397;
  assign or_690_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | or_tmp_398;
  assign or_685_nl = while_mux_1249_tmp | or_tmp_393;
  assign mux_tmp_296 = MUX_s_1_2_2(or_690_nl, or_685_nl, while_stage_0_5);
  assign mux_tmp_297 = MUX_s_1_2_2(or_tmp_398, or_tmp_393, while_stage_0_5);
  assign or_703_nl = weight_mem_read_arbxbar_arbiters_next_0_5_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]))
      | or_tmp_396;
  assign or_692_nl = weight_mem_read_arbxbar_arbiters_next_0_6_sva | or_tmp_397;
  assign mux_299_nl = MUX_s_1_2_2(or_703_nl, or_692_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign or_704_nl = while_mux_1251_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]))
      | or_tmp_391;
  assign or_691_nl = while_mux_1250_tmp | or_tmp_392;
  assign mux_298_nl = MUX_s_1_2_2(or_704_nl, or_691_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign mux_300_nl = MUX_s_1_2_2(mux_299_nl, mux_298_nl, while_stage_0_5);
  assign mux_301_nl = MUX_s_1_2_2(mux_300_nl, mux_tmp_297, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign mux_302_nl = MUX_s_1_2_2(mux_301_nl, mux_tmp_296, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign and_dcpl_648 = ~(mux_302_nl | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp);
  assign mux_303_nl = MUX_s_1_2_2(or_tmp_396, or_tmp_391, while_stage_0_5);
  assign and_dcpl_652 = (~ mux_303_nl) & (~(weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0])))
      & nor_253_cse;
  assign and_dcpl_655 = weight_mem_read_arbxbar_xbar_1_for_3_2_operator_7_false_1_operator_7_false_1_or_tmp
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_tmp);
  assign and_dcpl_656 = (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_7_false_1_operator_7_false_1_or_tmp)
      & weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_tmp;
  assign and_dcpl_657 = ~(weight_mem_read_arbxbar_xbar_1_for_3_2_operator_7_false_1_operator_7_false_1_or_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_tmp);
  assign and_dcpl_661 = (~(weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp))
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_3_Arbiter_8U_Roundrobin_pick_1_priority_and_6_tmp)
      & weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp;
  assign and_dcpl_662 = ~((~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]))) | weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp);
  assign and_dcpl_665 = nor_246_cse & (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]))
      & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp));
  assign or_dcpl_296 = ~(Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs);
  assign PECore_PushAxiRsp_mux_13_itm_1_mx0c1 = (~ rva_in_reg_rw_sva_5) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_a = weight_port_read_out_data_3_7_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[63:56];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_c = weight_port_read_out_data_3_6_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[55:48];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_1_a = weight_port_read_out_data_7_1_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[15:8];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_1_c = weight_port_read_out_data_7_0_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[7:0];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_2_a = weight_port_read_out_data_7_3_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[31:24];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_2_c = weight_port_read_out_data_7_2_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[23:16];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_3_a = weight_port_read_out_data_7_5_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[47:40];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_3_c = weight_port_read_out_data_7_4_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[39:32];
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_4_a = weight_port_read_out_data_7_7_sva_dfm_2;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_4_c = weight_port_read_out_data_7_6_sva_dfm_2;
  assign weight_port_read_out_data_mux_48_nl = MUX_s_1_2_2(weight_port_read_out_data_0_1_sva_dfm_2_7,
      Datapath_for_4_ProductSum_for_acc_5_cmp_5_a_mx1_7, fsm_output);
  assign weight_port_read_out_data_mux_75_nl = MUX_v_7_2_2(weight_port_read_out_data_0_1_sva_dfm_2_6_0,
      Datapath_for_4_ProductSum_for_acc_5_cmp_5_a_mx1_6_0, fsm_output);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_5_a = {weight_port_read_out_data_mux_48_nl
      , weight_port_read_out_data_mux_75_nl};
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_5_c = {weight_port_read_out_data_0_0_sva_dfm_3_7
      , weight_port_read_out_data_0_0_sva_dfm_3_6_0};
  assign weight_port_read_out_data_mux_47_nl = MUX_s_1_2_2(weight_port_read_out_data_0_3_sva_dfm_2_7_1,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_7, fsm_output);
  assign weight_port_read_out_data_mux_76_nl = MUX_v_3_2_2(weight_port_read_out_data_0_3_sva_dfm_2_6_4,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_6_4, fsm_output);
  assign weight_port_read_out_data_mux_77_nl = MUX_v_4_2_2(weight_port_read_out_data_0_3_sva_dfm_2_3_0,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_3_0, fsm_output);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_a = {weight_port_read_out_data_mux_47_nl
      , weight_port_read_out_data_mux_76_nl , weight_port_read_out_data_mux_77_nl};
  assign weight_port_read_out_data_mux_46_nl = MUX_s_1_2_2(weight_port_read_out_data_0_2_sva_dfm_2_7_1,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_7, fsm_output);
  assign weight_port_read_out_data_mux_78_nl = MUX_s_1_2_2(weight_port_read_out_data_0_2_sva_dfm_2_6,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_6, fsm_output);
  assign weight_port_read_out_data_mux_79_nl = MUX_v_6_2_2(weight_port_read_out_data_0_2_sva_dfm_2_5_0,
      Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_5_0, fsm_output);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_c = {weight_port_read_out_data_mux_46_nl
      , weight_port_read_out_data_mux_78_nl , weight_port_read_out_data_mux_79_nl};
  assign weight_port_read_out_data_mux_45_nl = MUX_v_4_2_2(weight_port_read_out_data_0_5_sva_dfm_2_7_4,
      Datapath_for_4_ProductSum_for_acc_5_cmp_7_a_mx1_7_4, fsm_output);
  assign weight_port_read_out_data_mux_80_nl = MUX_v_4_2_2(weight_port_read_out_data_0_5_sva_dfm_2_3_0,
      Datapath_for_4_ProductSum_for_acc_5_cmp_7_a_mx1_3_0, fsm_output);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_a = {weight_port_read_out_data_mux_45_nl
      , weight_port_read_out_data_mux_80_nl};
  assign weight_port_read_out_data_mux_44_nl = MUX_s_1_2_2(weight_port_read_out_data_0_4_sva_dfm_2_7,
      Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_7, fsm_output);
  assign weight_port_read_out_data_mux_81_nl = MUX_s_1_2_2(weight_port_read_out_data_0_4_sva_dfm_2_6,
      Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_6, fsm_output);
  assign weight_port_read_out_data_mux_82_nl = MUX_v_6_2_2(weight_port_read_out_data_0_4_sva_dfm_2_5_0,
      Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_5_0, fsm_output);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_c = {weight_port_read_out_data_mux_44_nl
      , weight_port_read_out_data_mux_81_nl , weight_port_read_out_data_mux_82_nl};
  assign weight_port_read_out_data_mux_43_nl = MUX_s_1_2_2(weight_port_read_out_data_0_7_sva_dfm_2_7,
      Datapath_for_4_ProductSum_for_acc_5_cmp_8_a_mx1_7, fsm_output);
  assign weight_port_read_out_data_mux_83_nl = MUX_v_7_2_2(weight_port_read_out_data_0_7_sva_dfm_2_6_0,
      Datapath_for_4_ProductSum_for_acc_5_cmp_8_a_mx1_6_0, fsm_output);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_8_a = {weight_port_read_out_data_mux_43_nl
      , weight_port_read_out_data_mux_83_nl};
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_8_c = MUX_v_8_2_2(({weight_port_read_out_data_0_6_sva_dfm_2_7_4
      , weight_port_read_out_data_0_6_sva_dfm_2_3_0}), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000,
      weight_mem_run_3_for_land_1_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_9_a = MUX_v_8_2_2(weight_port_read_out_data_6_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_9_c = MUX_v_8_2_2(weight_port_read_out_data_6_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_10_a = MUX_v_8_2_2(weight_port_read_out_data_6_3_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_10_c = MUX_v_8_2_2(weight_port_read_out_data_6_2_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_11_a = MUX_v_8_2_2(weight_port_read_out_data_6_5_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_11_c = MUX_v_8_2_2(weight_port_read_out_data_6_4_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_12_a = MUX_v_8_2_2(weight_port_read_out_data_6_7_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_12_c = MUX_v_8_2_2(weight_port_read_out_data_6_6_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_13_a = MUX_v_8_2_2(weight_port_read_out_data_1_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_13_c = MUX_v_8_2_2(weight_port_read_out_data_1_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_14_a = MUX_v_8_2_2(weight_port_read_out_data_1_3_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_14_c = MUX_v_8_2_2(weight_port_read_out_data_1_2_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_15_a = MUX_v_8_2_2(weight_port_read_out_data_1_5_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_15_c = MUX_v_8_2_2(weight_port_read_out_data_1_4_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_16_a = MUX_v_8_2_2(weight_port_read_out_data_1_7_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_000000,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_16_c = MUX_v_8_2_2(weight_port_read_out_data_1_6_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_17_a = weight_port_read_out_data_5_1_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_17_c = weight_port_read_out_data_5_0_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_18_a = weight_port_read_out_data_5_3_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_18_c = weight_port_read_out_data_5_2_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_19_a = weight_port_read_out_data_5_5_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_19_c = weight_port_read_out_data_5_4_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_20_a = weight_port_read_out_data_5_7_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_20_c = weight_port_read_out_data_5_6_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_21_a = {weight_mem_run_3_for_5_mux_17_itm_1_7
      , weight_mem_run_3_for_5_mux_17_itm_1_6 , weight_mem_run_3_for_5_mux_17_itm_1_5_0};
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_21_b = {input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_7
      , input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_6_0};
  assign and_527_nl = fsm_output & (~ weight_mem_run_3_for_land_3_lpi_1_dfm_3);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_21_c = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000,
      weight_port_read_out_data_2_0_sva_dfm_1, and_527_nl);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_21_d = {input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_7
      , input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_6_0};
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_22_a = MUX_v_8_2_2(weight_port_read_out_data_2_3_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001,
      weight_mem_run_3_for_land_3_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_22_c = MUX_v_8_2_2(weight_port_read_out_data_2_2_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002,
      weight_mem_run_3_for_land_3_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_23_a = MUX_v_8_2_2(weight_port_read_out_data_2_5_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003,
      weight_mem_run_3_for_land_3_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_23_c = MUX_v_8_2_2(weight_port_read_out_data_2_4_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004,
      weight_mem_run_3_for_land_3_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_24_a = MUX_v_8_2_2(weight_port_read_out_data_2_7_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_sva_1,
      weight_mem_run_3_for_land_3_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_24_c = MUX_v_8_2_2(weight_port_read_out_data_2_6_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005,
      weight_mem_run_3_for_land_3_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_25_a = MUX_v_8_2_2(weight_port_read_out_data_4_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_25_c = MUX_v_8_2_2(weight_port_read_out_data_4_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_26_a = MUX_v_8_2_2(weight_port_read_out_data_4_3_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_26_c = MUX_v_8_2_2(weight_port_read_out_data_4_2_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_27_a = MUX_v_8_2_2(weight_port_read_out_data_4_5_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_27_c = MUX_v_8_2_2(weight_port_read_out_data_4_4_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_28_a = MUX_v_8_2_2(weight_port_read_out_data_4_7_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_28_c = MUX_v_8_2_2(weight_port_read_out_data_4_6_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_29_a = MUX_v_8_2_2(weight_port_read_out_data_3_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_29_c = MUX_v_8_2_2(weight_port_read_out_data_3_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_30_a = MUX_v_8_2_2(weight_port_read_out_data_3_3_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_30_c = MUX_v_8_2_2(weight_port_read_out_data_3_2_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_31_a = weight_port_read_out_data_3_5_sva_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_31_c = weight_port_read_out_data_3_4_sva_dfm_3;
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0));
  assign weight_mem_banks_write_if_for_if_and_35_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_36_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_37_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_38_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_39_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_40_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_41_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      , weight_mem_banks_write_if_for_if_and_35_nl , weight_mem_banks_write_if_for_if_and_36_nl
      , weight_mem_banks_write_if_for_if_and_37_nl , weight_mem_banks_write_if_for_if_and_38_nl
      , weight_mem_banks_write_if_for_if_and_39_nl , weight_mem_banks_write_if_for_if_and_40_nl
      , weight_mem_banks_write_if_for_if_and_41_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0});
  assign weight_mem_banks_write_if_for_if_mux_7_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      , weight_mem_banks_write_if_for_if_mux_7_nl};
  assign nor_412_nl = ~((~ PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3) |
      PECore_RunFSM_switch_lp_equal_tmp_1_2);
  assign mux_151_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse,
      nor_412_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff = mux_151_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_2[14:3];
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff = and_dcpl_170;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0));
  assign weight_mem_banks_write_if_for_if_and_28_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_29_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_30_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_31_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_32_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_33_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_34_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      , weight_mem_banks_write_if_for_if_and_28_nl , weight_mem_banks_write_if_for_if_and_29_nl
      , weight_mem_banks_write_if_for_if_and_30_nl , weight_mem_banks_write_if_for_if_and_31_nl
      , weight_mem_banks_write_if_for_if_and_32_nl , weight_mem_banks_write_if_for_if_and_33_nl
      , weight_mem_banks_write_if_for_if_and_34_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0});
  assign weight_mem_banks_write_if_for_if_mux_6_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      , weight_mem_banks_write_if_for_if_mux_6_nl};
  assign nor_411_nl = ~(PECore_UpdateFSM_switch_lp_equal_tmp_2_3 | (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_150_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse,
      nor_411_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff = mux_150_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff = and_dcpl_173;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0));
  assign weight_mem_banks_write_if_for_if_and_21_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_22_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_23_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_24_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_25_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_26_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_27_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      , weight_mem_banks_write_if_for_if_and_21_nl , weight_mem_banks_write_if_for_if_and_22_nl
      , weight_mem_banks_write_if_for_if_and_23_nl , weight_mem_banks_write_if_for_if_and_24_nl
      , weight_mem_banks_write_if_for_if_and_25_nl , weight_mem_banks_write_if_for_if_and_26_nl
      , weight_mem_banks_write_if_for_if_and_27_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0});
  assign weight_mem_banks_write_if_for_if_mux_5_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      , weight_mem_banks_write_if_for_if_mux_5_nl};
  assign nor_410_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_3) | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]));
  assign mux_149_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse,
      nor_410_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff = mux_149_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff = and_dcpl_176;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0));
  assign weight_mem_banks_write_if_for_if_and_14_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_15_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_16_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_17_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_18_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_19_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_20_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      , weight_mem_banks_write_if_for_if_and_14_nl , weight_mem_banks_write_if_for_if_and_15_nl
      , weight_mem_banks_write_if_for_if_and_16_nl , weight_mem_banks_write_if_for_if_and_17_nl
      , weight_mem_banks_write_if_for_if_and_18_nl , weight_mem_banks_write_if_for_if_and_19_nl
      , weight_mem_banks_write_if_for_if_and_20_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0});
  assign weight_mem_banks_write_if_for_if_mux_4_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      , weight_mem_banks_write_if_for_if_mux_4_nl};
  assign nor_409_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3) | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]));
  assign mux_148_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse,
      nor_409_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff = mux_148_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff = and_dcpl_179;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0));
  assign weight_mem_banks_write_if_for_if_and_7_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_9_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_10_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_11_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_12_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_13_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      , weight_mem_banks_write_if_for_if_and_7_nl , weight_mem_banks_write_if_for_if_and_8_nl
      , weight_mem_banks_write_if_for_if_and_9_nl , weight_mem_banks_write_if_for_if_and_10_nl
      , weight_mem_banks_write_if_for_if_and_11_nl , weight_mem_banks_write_if_for_if_and_12_nl
      , weight_mem_banks_write_if_for_if_and_13_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0});
  assign weight_mem_banks_write_if_for_if_mux_3_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      , weight_mem_banks_write_if_for_if_mux_3_nl};
  assign or_406_nl = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp;
  assign or_405_nl = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp;
  assign mux_146_nl = MUX_s_1_2_2(or_406_nl, or_405_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign or_710_nl = Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp | mux_146_nl;
  assign nor_408_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1)
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]));
  assign mux_147_nl = MUX_s_1_2_2(or_710_nl, nor_408_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff = mux_147_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff = and_dcpl_182;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0));
  assign weight_mem_banks_write_if_for_if_and_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_1_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_2_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_3_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_5_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl ,
      weight_mem_banks_write_if_for_if_and_nl , weight_mem_banks_write_if_for_if_and_1_nl
      , weight_mem_banks_write_if_for_if_and_2_nl , weight_mem_banks_write_if_for_if_and_3_nl
      , weight_mem_banks_write_if_for_if_and_4_nl , weight_mem_banks_write_if_for_if_and_5_nl
      , weight_mem_banks_write_if_for_if_and_6_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0});
  assign weight_mem_banks_write_if_for_if_mux_2_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      , weight_mem_banks_write_if_for_if_mux_2_nl};
  assign nor_406_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1)
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]));
  assign mux_145_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse,
      nor_406_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff = mux_145_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff = and_dcpl_185;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_1_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_54_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0,
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_1_nl
      , weight_mem_banks_write_if_for_if_mux_54_nl};
  assign nor_405_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1));
  assign mux_144_nl = MUX_s_1_2_2(mux_tmp_102, nor_405_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff = mux_144_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_3_14_3;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff = and_dcpl_489;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_53_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0,
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_nl
      , weight_mem_banks_write_if_for_if_mux_53_nl};
  assign nor_404_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1));
  assign mux_143_nl = MUX_s_1_2_2(mux_tmp_98, nor_404_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff = mux_143_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff = and_dcpl_486;
  assign or_dcpl_297 = ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]) & and_dcpl_594)
      | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]) & and_dcpl_597) | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[2])
      & and_dcpl_595);
  assign and_dcpl_678 = (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1;
  assign and_dcpl_679 = (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1;
  assign or_dcpl_302 = and_dcpl_679 | and_dcpl_678;
  assign or_dcpl_303 = and_dcpl_679 | ((pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1);
  assign PECore_DecodeAxiRead_switch_lp_mux_21_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[0]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl
      = PECore_DecodeAxiRead_switch_lp_mux_21_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_20_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl,
      rva_out_reg_data_0_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_14_itm = MUX_s_1_2_2(rva_out_reg_data_mux_20_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl
      = (SC_SRAM_CONFIG[7]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9) &
      PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_10_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl,
      rva_out_reg_data_7_1_sva_dfm_6_6, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3[6]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_6, {PECore_PushAxiRsp_if_asn_55
      , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl
      = (SC_SRAM_CONFIG[6:1]) & (signext_6_1(~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9))
      & ({{5{PECore_DecodeAxiRead_switch_lp_nor_9_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1});
  assign PECore_PushAxiRsp_if_mux1h_10_5_0 = MUX1HOT_v_6_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl,
      rva_out_reg_data_7_1_sva_dfm_6_5_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3[5:0]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_5_0,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_22_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[8]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl
      = PECore_DecodeAxiRead_switch_lp_mux_22_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_21_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl,
      rva_out_reg_data_8_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_15_itm = MUX_s_1_2_2(rva_out_reg_data_mux_21_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_DecodeAxiRead_switch_lp_mux_18_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[15]),
      rva_out_reg_data_15_9_sva_dfm_10_6, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl
      = PECore_DecodeAxiRead_switch_lp_mux_18_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_12_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl,
      rva_out_reg_data_15_9_sva_dfm_6_6, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3[6]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_6, {PECore_PushAxiRsp_if_asn_55
      , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_26_nl = MUX_v_6_2_2((SC_SRAM_CONFIG[14:9]),
      rva_out_reg_data_15_9_sva_dfm_10_5_0, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl
      = MUX_v_6_2_2(6'b000000, PECore_DecodeAxiRead_switch_lp_mux_26_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_12_5_0 = MUX1HOT_v_6_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl,
      rva_out_reg_data_15_9_sva_dfm_6_5_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3[5:0]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_5_0,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_23_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[16]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl
      = PECore_DecodeAxiRead_switch_lp_mux_23_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_22_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl,
      rva_out_reg_data_16_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_16_itm = MUX_s_1_2_2(rva_out_reg_data_mux_22_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_DecodeAxiRead_switch_lp_mux_24_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[24]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl
      = PECore_DecodeAxiRead_switch_lp_mux_24_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_24_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl,
      rva_out_reg_data_24_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_17_nl = MUX_s_1_2_2(rva_out_reg_data_mux_24_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_PushAxiRsp_if_mux1h_15 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_17_nl,
      (weight_port_read_out_data_0_3_sva_dfm_5_6_0_rsp_1[0]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign PECore_DecodeAxiRead_switch_lp_mux_20_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[30:28]),
      (rva_out_reg_data_30_25_sva_dfm_8[5:3]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl =
      MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_20_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_16_5_3 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl,
      rva_out_reg_data_30_25_sva_dfm_6_5_3, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3[5:3]),
      weight_port_read_out_data_0_3_sva_dfm_5_6_0_rsp_0, {PECore_PushAxiRsp_if_asn_55
      , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_27_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[27:25]),
      (rva_out_reg_data_30_25_sva_dfm_8[2:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl
      = MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_27_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_16_2_0 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl,
      rva_out_reg_data_30_25_sva_dfm_6_2_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3[2:0]),
      (weight_port_read_out_data_0_3_sva_dfm_5_6_0_rsp_1[3:1]), {PECore_PushAxiRsp_if_asn_55
      , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl
      = (SC_SRAM_CONFIG[31]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9) &
      PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_23_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl,
      rva_out_reg_data_31_sva_dfm_6, rva_in_reg_rw_sva_10);
  assign PECore_PushAxiRsp_if_else_mux_18_nl = MUX_s_1_2_2(rva_out_reg_data_mux_23_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3,
      input_read_req_valid_lpi_1_dfm_1_10);
  assign PECore_PushAxiRsp_if_mux1h_17 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_18_nl,
      weight_port_read_out_data_0_3_sva_dfm_5_7, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
  assign or_5_nl = rva_in_reg_rw_sva_st_1_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5
      | rva_in_reg_rw_sva_5 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1;
  assign mux_2_nl = MUX_s_1_2_2((~ PECore_RunMac_PECore_RunMac_if_and_svs_st_5),
      or_5_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_3_nl = MUX_s_1_2_2(or_tmp, mux_2_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4);
  assign mux_4_nl = MUX_s_1_2_2(mux_3_nl, mux_tmp, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign weight_mem_run_3_for_5_and_222_ssc = PECoreRun_wen & (~ mux_4_nl) & while_stage_0_7;
  assign mux_58_nl = MUX_s_1_2_2((~ or_tmp_84), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign weight_mem_banks_load_store_for_else_and_1_ssc = PECoreRun_wen & mux_58_nl
      & and_dcpl_43;
  assign mux_61_nl = MUX_s_1_2_2(or_tmp_84, mux_tmp_60, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign weight_mem_banks_load_store_for_else_and_7_ssc = PECoreRun_wen & (~ mux_61_nl)
      & and_dcpl_43;
  assign or_241_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1 |
      rva_in_reg_rw_sva_st_1_4 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4
      | (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3) | PECore_DecodeAxiRead_switch_lp_nor_tmp_4
      | rva_in_reg_rw_sva_4;
  assign mux_69_nl = MUX_s_1_2_2(or_241_nl, mux_tmp_60, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign weight_mem_banks_load_store_for_else_and_17_ssc = PECoreRun_wen & (~ mux_69_nl)
      & and_dcpl_43;
  assign weight_port_read_out_data_and_94_ssc = PECoreRun_wen & ((and_dcpl_350 &
      (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 | PECore_DecodeAxiRead_switch_lp_nor_tmp_5))
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 | rva_in_reg_rw_sva_st_1_5))
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4) | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      & and_dcpl_357;
  assign mux1h_nl = MUX1HOT_s_1_8_2((rva_out_reg_data_55_48_sva_dfm_1_5[7]), (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[15]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[15]),
      weight_port_read_out_data_0_1_sva_dfm_2_7, {and_927_cse , and_928_cse , and_929_cse
      , and_930_cse , and_931_cse , and_932_cse , and_933_cse , nor_426_cse});
  assign weight_port_read_out_data_0_1_sva_dfm_mx0w1_7 = mux1h_nl & (~ or_dcpl_302);
  assign mux1h_8_nl = MUX1HOT_v_7_8_2((rva_out_reg_data_55_48_sva_dfm_1_5[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[14:8]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[14:8]),
      weight_port_read_out_data_0_1_sva_dfm_2_6_0, {and_927_cse , and_928_cse , and_929_cse
      , and_930_cse , and_931_cse , and_932_cse , and_933_cse , nor_426_cse});
  assign not_2301_nl = ~ or_dcpl_302;
  assign weight_port_read_out_data_0_1_sva_dfm_mx0w1_6_0 = MUX_v_7_2_2(7'b0000000,
      mux1h_8_nl, not_2301_nl);
  assign and_936_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 & (~ or_dcpl_303);
  assign mux1h_2_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[7]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[7]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[7]),
      weight_port_read_out_data_0_0_sva_dfm_2_7, {and_936_ssc , and_937_cse , and_938_cse
      , and_939_cse , and_940_cse , and_941_cse , and_942_cse , nor_427_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w1_7 = mux1h_2_nl & (~ or_dcpl_303);
  assign mux1h_9_nl = MUX1HOT_v_7_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[6:0]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[6:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[6:0]),
      weight_port_read_out_data_0_0_sva_dfm_2_6_0, {and_936_ssc , and_937_cse , and_938_cse
      , and_939_cse , and_940_cse , and_941_cse , and_942_cse , nor_427_cse});
  assign not_2302_nl = ~ or_dcpl_303;
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w1_6_0 = MUX_v_7_2_2(7'b0000000,
      mux1h_9_nl, not_2302_nl);
  assign and_945_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_dcpl_303);
  assign mux1h_3_nl = MUX1HOT_s_1_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6[1]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[23]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[23]),
      weight_port_read_out_data_0_2_sva_dfm_2_7_1, {and_945_ssc , and_937_cse , and_938_cse
      , and_939_cse , and_940_cse , and_941_cse , and_942_cse , nor_427_cse});
  assign weight_port_read_out_data_0_2_sva_dfm_mx0w2_7 = mux1h_3_nl & (~ or_dcpl_303);
  assign mux1h_10_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6[0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[6]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[22]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[22]),
      weight_port_read_out_data_0_2_sva_dfm_2_6, {and_945_ssc , and_937_cse , and_938_cse
      , and_939_cse , and_940_cse , and_941_cse , and_942_cse , nor_427_cse});
  assign weight_port_read_out_data_0_2_sva_dfm_mx0w2_6 = mux1h_10_nl & (~ or_dcpl_303);
  assign mux1h_11_nl = MUX1HOT_v_6_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0[5:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[5:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[21:16]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[21:16]),
      weight_port_read_out_data_0_2_sva_dfm_2_5_0, {and_945_ssc , and_937_cse , and_938_cse
      , and_939_cse , and_940_cse , and_941_cse , and_942_cse , nor_427_cse});
  assign not_2303_nl = ~ or_dcpl_303;
  assign weight_port_read_out_data_0_2_sva_dfm_mx0w2_5_0 = MUX_v_6_2_2(6'b000000,
      mux1h_11_nl, not_2303_nl);
  assign mux1h_4_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4[3]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[31]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[31]),
      weight_port_read_out_data_0_3_sva_dfm_2_7_1, {and_927_cse , and_928_cse , and_929_cse
      , and_930_cse , and_931_cse , and_932_cse , and_933_cse , nor_426_cse});
  assign weight_port_read_out_data_0_3_sva_dfm_mx0w0_7 = mux1h_4_nl & (~ or_dcpl_302);
  assign mux1h_12_nl = MUX1HOT_v_3_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[6:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0[6:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4[2:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[6:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[6:4]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[30:28]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[30:28]),
      weight_port_read_out_data_0_3_sva_dfm_2_6_4, {and_927_cse , and_928_cse , and_929_cse
      , and_930_cse , and_931_cse , and_932_cse , and_933_cse , nor_426_cse});
  assign not_2305_nl = ~ or_dcpl_302;
  assign weight_port_read_out_data_0_3_sva_dfm_mx0w0_6_4 = MUX_v_3_2_2(3'b000, mux1h_12_nl,
      not_2305_nl);
  assign mux1h_13_nl = MUX1HOT_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[3:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[27:24]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[27:24]),
      weight_port_read_out_data_0_3_sva_dfm_2_3_0, {and_927_cse , and_928_cse , and_929_cse
      , and_930_cse , and_931_cse , and_932_cse , and_933_cse , nor_426_cse});
  assign not_2306_nl = ~ or_dcpl_302;
  assign weight_port_read_out_data_0_3_sva_dfm_mx0w0_3_0 = MUX_v_4_2_2(4'b0000, mux1h_13_nl,
      not_2306_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_136_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[55:52]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_136_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_137_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[55:52]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_137_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_7_4
      = MUX_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7_4,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_87_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_64_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[51:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_87_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_80_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_65_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[51:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_80_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_3_0
      = MUX_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_64_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_65_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign mux1h_5_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[63]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63]),
      weight_port_read_out_data_0_7_sva_dfm_2_7, {and_927_cse , and_928_cse , and_929_cse
      , and_930_cse , and_931_cse , and_932_cse , and_933_cse , nor_426_cse});
  assign weight_port_read_out_data_0_7_sva_dfm_3_7 = mux1h_5_nl & (~ or_dcpl_302);
  assign mux1h_14_nl = MUX1HOT_v_7_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[62:56]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[62:56]),
      weight_port_read_out_data_0_7_sva_dfm_2_6_0, {and_927_cse , and_928_cse , and_929_cse
      , and_930_cse , and_931_cse , and_932_cse , and_933_cse , nor_426_cse});
  assign not_2307_nl = ~ or_dcpl_302;
  assign weight_port_read_out_data_0_7_sva_dfm_3_6_0 = MUX_v_7_2_2(7'b0000000, mux1h_14_nl,
      not_2307_nl);
  assign and_972_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_718_tmp);
  assign and_973_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56 & (~ or_718_tmp);
  assign and_974_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse & (~ or_718_tmp);
  assign and_975_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      & (~ or_718_tmp);
  assign and_976_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1
      & (~ or_718_tmp);
  assign and_977_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1
      & (~ or_718_tmp);
  assign and_978_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      & (~ or_718_tmp);
  assign nor_431_ssc = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_718_tmp);
  assign mux1h_6_nl = MUX1HOT_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1[7:4]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[47:44]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[47:44]),
      weight_port_read_out_data_0_5_sva_dfm_2_7_4, {and_972_ssc , and_973_ssc , and_974_ssc
      , and_975_ssc , and_976_ssc , and_977_ssc , and_978_ssc , nor_431_ssc});
  assign not_2308_nl = ~ or_718_tmp;
  assign weight_port_read_out_data_0_5_sva_dfm_3_7_4 = MUX_v_4_2_2(4'b0000, mux1h_6_nl,
      not_2308_nl);
  assign mux1h_15_nl = MUX1HOT_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1[3:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[43:40]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[43:40]),
      weight_port_read_out_data_0_5_sva_dfm_2_3_0, {and_972_ssc , and_973_ssc , and_974_ssc
      , and_975_ssc , and_976_ssc , and_977_ssc , and_978_ssc , nor_431_ssc});
  assign not_2230_nl = ~ or_718_tmp;
  assign weight_port_read_out_data_0_5_sva_dfm_3_3_0 = MUX_v_4_2_2(4'b0000, mux1h_15_nl,
      not_2230_nl);
  assign and_981_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 & (~ or_dcpl_302);
  assign and_984_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      & (~ or_dcpl_302);
  assign and_985_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1
      & (~ or_dcpl_302);
  assign mux1h_7_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6[1]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[39]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[39]),
      weight_port_read_out_data_0_4_sva_dfm_2_7, {and_981_ssc , and_928_cse , and_929_cse
      , and_984_ssc , and_985_ssc , and_932_cse , and_933_cse , nor_426_cse});
  assign weight_port_read_out_data_0_4_sva_dfm_3_7 = mux1h_7_nl & (~ or_dcpl_302);
  assign mux1h_16_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6[0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1[6]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[38]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[38]),
      weight_port_read_out_data_0_4_sva_dfm_2_6, {and_981_ssc , and_928_cse , and_929_cse
      , and_984_ssc , and_985_ssc , and_932_cse , and_933_cse , nor_426_cse});
  assign weight_port_read_out_data_0_4_sva_dfm_3_6 = mux1h_16_nl & (~ or_dcpl_302);
  assign mux1h_17_nl = MUX1HOT_v_6_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[5:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1[5:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[37:32]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[37:32]),
      weight_port_read_out_data_0_4_sva_dfm_2_5_0, {and_981_ssc , and_928_cse , and_929_cse
      , and_984_ssc , and_985_ssc , and_932_cse , and_933_cse , nor_426_cse});
  assign not_2309_nl = ~ or_dcpl_302;
  assign weight_port_read_out_data_0_4_sva_dfm_3_5_0 = MUX_v_6_2_2(6'b000000, mux1h_17_nl,
      not_2309_nl);
  assign mux_1_nl = MUX_s_1_2_2(or_tmp, mux_tmp, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign input_mem_banks_read_1_read_data_and_ssc = PECoreRun_wen & (~ mux_1_nl)
      & while_stage_0_7;
  assign weight_port_read_out_data_and_1_ssc = PECoreRun_wen & ((weight_mem_run_3_for_land_1_lpi_1_dfm_3
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5))
      | while_and_24_cse) & while_stage_0_7;
  assign or_2319_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1;
  assign or_2318_nl = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1;
  assign mux_885_nl = MUX_s_1_2_2(or_2319_nl, or_2318_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign or_2317_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse |
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1;
  assign mux_886_nl = MUX_s_1_2_2(mux_885_nl, or_2317_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign and_1831_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & mux_886_nl;
  assign or_2320_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1 | and_1831_cse;
  assign and_2186_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2
      | reg_weight_mem_run_3_for_5_and_167_itm_2_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign or_2327_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1 | and_1831_cse;
  assign mux_890_nl = MUX_s_1_2_2(and_2186_nl, or_2327_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_1835_cse = mux_890_nl & weight_mem_run_3_for_aelse_and_cse;
  assign or_2340_nl = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1;
  assign or_2339_nl = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1;
  assign mux_894_nl = MUX_s_1_2_2(or_2340_nl, or_2339_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign or_2338_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse |
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1;
  assign mux_895_nl = MUX_s_1_2_2(mux_894_nl, or_2338_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign and_1840_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & mux_895_nl;
  assign and_2190_cse = (reg_weight_mem_run_3_for_5_and_168_itm_2_cse | reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_166_itm_2_cse | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_162_itm_2_cse | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_port_read_out_data_and_99_enex5 = weight_port_read_out_data_and_86_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo;
  assign weight_port_read_out_data_and_100_enex5 = weight_port_read_out_data_and_86_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo;
  assign rva_out_reg_data_and_126_enex5 = rva_out_reg_data_and_34_cse & reg_rva_out_reg_data_23_17_sva_dfm_5_1_enexo;
  assign rva_out_reg_data_and_127_enex5 = rva_out_reg_data_and_34_cse & reg_rva_out_reg_data_15_9_sva_dfm_7_1_enexo;
  assign rva_out_reg_data_and_128_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_129_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_130_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_131_enex5 = rva_out_reg_data_and_42_cse & reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_132_enex5 = rva_out_reg_data_and_42_cse & reg_weight_mem_run_3_for_5_mux_17_itm_1_2_enexo;
  assign weight_port_read_out_data_and_90_ssc = PECoreRun_wen & and_dcpl_30 & (~
      rva_in_reg_rw_sva_st_1_6) & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
  assign weight_port_read_out_data_and_101_enex5 = weight_port_read_out_data_and_90_ssc
      & reg_input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_1_enexo;
  assign weight_port_read_out_data_and_102_enex5 = weight_port_read_out_data_and_90_ssc
      & reg_input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_1_enexo;
  assign rva_out_reg_data_and_133_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_1_1_enexo;
  assign rva_out_reg_data_and_134_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_135_enex5 = input_read_req_valid_and_3_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_1_1_enexo;
  assign weight_mem_run_3_for_5_and_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_179_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_180_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_181_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_8_a_mx1_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_7_sva_dfm_2_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_ssc
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_179_ssc
      , weight_mem_run_3_for_5_and_180_ssc , weight_mem_run_3_for_5_and_181_ssc});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_8_a_mx1_6_0 = MUX1HOT_v_7_9_2(weight_port_read_out_data_0_7_sva_dfm_2_6_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[62:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[62:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[62:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[62:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[62:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[62:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[62:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[54:48]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_ssc
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_179_ssc
      , weight_mem_run_3_for_5_and_180_ssc , weight_mem_run_3_for_5_and_181_ssc});
  assign weight_mem_run_3_for_5_and_187_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_188_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_4_sva_dfm_2_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[39]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_187_ssc
      , weight_mem_run_3_for_5_and_188_ssc , weight_mem_run_3_for_5_and_189_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_6 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_4_sva_dfm_2_6,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[38]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[38]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[38]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[38]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[38]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[38]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[38]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[30]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_187_ssc
      , weight_mem_run_3_for_5_and_188_ssc , weight_mem_run_3_for_5_and_189_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_5_0 = MUX1HOT_v_6_9_2(weight_port_read_out_data_0_4_sva_dfm_2_5_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[37:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[37:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[37:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[37:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[37:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[37:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[37:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[29:24]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_187_ssc
      , weight_mem_run_3_for_5_and_188_ssc , weight_mem_run_3_for_5_and_189_cse});
  assign weight_mem_run_3_for_5_and_190_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_191_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_192_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_193_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_194_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_195_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_a_mx1_7_4 = MUX1HOT_v_4_9_2(weight_port_read_out_data_0_5_sva_dfm_2_7_4,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:44]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:44]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:44]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:44]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:44]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:44]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:44]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:36]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_190_ssc
      , weight_mem_run_3_for_5_and_191_ssc , weight_mem_run_3_for_5_and_192_ssc ,
      weight_mem_run_3_for_5_and_193_ssc , weight_mem_run_3_for_5_and_194_ssc , weight_mem_run_3_for_5_and_195_ssc
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_197_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_7_a_mx1_3_0 = MUX1HOT_v_4_9_2(weight_port_read_out_data_0_5_sva_dfm_2_3_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[43:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[43:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[43:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[43:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[43:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[43:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[43:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[35:32]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_190_ssc
      , weight_mem_run_3_for_5_and_191_ssc , weight_mem_run_3_for_5_and_192_ssc ,
      weight_mem_run_3_for_5_and_193_ssc , weight_mem_run_3_for_5_and_194_ssc , weight_mem_run_3_for_5_and_195_ssc
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_197_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_2_sva_dfm_2_7_1,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[23]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_203_cse
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_189_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_6 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_2_sva_dfm_2_6,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[22]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[22]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[22]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[22]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[22]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[22]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[22]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[14]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_203_cse
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_189_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_5_0 = MUX1HOT_v_6_9_2(weight_port_read_out_data_0_2_sva_dfm_2_5_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[21:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[21:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[21:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[21:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[21:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[21:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[21:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[13:8]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_203_cse
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_189_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_3_sva_dfm_2_7_1,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[31]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_203_cse
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_197_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_6_4 = MUX1HOT_v_3_9_2(weight_port_read_out_data_0_3_sva_dfm_2_6_4,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[30:28]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[30:28]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[30:28]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[30:28]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[30:28]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[30:28]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[30:28]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[22:20]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_203_cse
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_197_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_3_0 = MUX1HOT_v_4_9_2(weight_port_read_out_data_0_3_sva_dfm_2_3_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[27:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[27:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[27:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[27:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[27:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[27:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[27:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[19:16]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_203_cse
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_197_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_3_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_0_sva_dfm_2_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[7]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[7]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , reg_weight_mem_run_3_for_5_and_162_itm_2_cse , reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      , weight_mem_run_3_for_5_and_164_itm_2 , reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_166_itm_2_cse , reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_168_itm_2_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_3_6_0 = MUX1HOT_v_7_9_2(weight_port_read_out_data_0_0_sva_dfm_2_6_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[6:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[6:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[6:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[6:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[6:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[6:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[6:0]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[6:0]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , reg_weight_mem_run_3_for_5_and_162_itm_2_cse , reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      , weight_mem_run_3_for_5_and_164_itm_2 , reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_166_itm_2_cse , reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_168_itm_2_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_5_a_mx1_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_1_sva_dfm_2_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[15]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_203_cse
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_189_cse});
  assign Datapath_for_4_ProductSum_for_acc_5_cmp_5_a_mx1_6_0 = MUX1HOT_v_7_9_2(weight_port_read_out_data_0_1_sva_dfm_2_6_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[14:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[14:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[14:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[14:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[14:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[14:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[14:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[6:0]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_203_cse
      , weight_mem_run_3_for_5_and_196_cse , weight_mem_run_3_for_5_and_189_cse});
  assign rva_out_reg_data_55_48_sva_dfm_6_mx1_7_4 = MUX_v_4_2_2(rva_out_reg_data_55_48_sva_dfm_4_1_7_4,
      rva_out_reg_data_55_48_sva_dfm_6_rsp_0, or_dcpl_283);
  assign rva_out_reg_data_55_48_sva_dfm_6_mx1_3_0 = MUX_v_4_2_2(rva_out_reg_data_55_48_sva_dfm_4_1_3_0,
      rva_out_reg_data_55_48_sva_dfm_6_rsp_1, or_dcpl_283);
  assign rva_out_reg_data_46_40_sva_dfm_6_mx1_6_4 = MUX_v_3_2_2(rva_out_reg_data_46_40_sva_dfm_4_1_6_4,
      rva_out_reg_data_46_40_sva_dfm_6_rsp_0, or_dcpl_283);
  assign rva_out_reg_data_46_40_sva_dfm_6_mx1_3_0 = MUX_v_4_2_2(rva_out_reg_data_46_40_sva_dfm_4_1_3_0,
      rva_out_reg_data_46_40_sva_dfm_6_rsp_1, or_dcpl_283);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1_3 = MUX_s_1_2_2(rva_out_reg_data_39_36_sva_dfm_4_1_3,
      rva_out_reg_data_39_36_sva_dfm_6_rsp_0, or_dcpl_283);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1_2 = MUX_s_1_2_2(rva_out_reg_data_39_36_sva_dfm_4_1_2,
      rva_out_reg_data_39_36_sva_dfm_6_rsp_1, or_dcpl_283);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1_1_0 = MUX_v_2_2_2(rva_out_reg_data_39_36_sva_dfm_4_1_1_0,
      rva_out_reg_data_39_36_sva_dfm_6_rsp_2, or_dcpl_283);
  assign weight_port_read_out_data_and_103_enex5 = weight_port_read_out_data_and_86_cse
      & reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo;
  assign weight_port_read_out_data_and_104_enex5 = weight_port_read_out_data_and_86_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_2_2_enexo;
  assign weight_port_read_out_data_and_105_enex5 = weight_port_read_out_data_and_90_ssc
      & reg_weight_mem_run_3_for_5_mux_17_itm_1_2_enexo_1;
  assign weight_port_read_out_data_and_106_enex5 = weight_port_read_out_data_and_90_ssc
      & reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo_1;
  assign rva_out_reg_data_and_136_enex5 = rva_out_reg_data_and_14_cse & reg_rva_out_reg_data_15_9_sva_dfm_9_1_enexo;
  assign rva_out_reg_data_and_137_enex5 = rva_out_reg_data_and_14_cse & reg_rva_out_reg_data_23_17_sva_dfm_7_1_enexo;
  assign rva_out_reg_data_and_138_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_4_enexo;
  assign rva_out_reg_data_and_139_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_4_1_enexo;
  assign rva_out_reg_data_and_140_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_4_1_enexo;
  assign weight_port_read_out_data_and_107_enex5 = weight_port_read_out_data_and_64_cse
      & reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_1_enexo;
  assign weight_port_read_out_data_and_108_enex5 = weight_port_read_out_data_and_64_cse
      & reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_1_enexo;
  assign PECore_DecodeAxiRead_switch_lp_mux_19_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[23]),
      (rva_out_reg_data_23_17_sva_dfm_8_6_4[2]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl
      = PECore_DecodeAxiRead_switch_lp_mux_19_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_14_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl,
      rva_out_reg_data_23_17_sva_dfm_6_6, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3[6]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_6, {PECore_PushAxiRsp_if_asn_55
      , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_25_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[22]),
      (rva_out_reg_data_23_17_sva_dfm_8_6_4[1]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl
      = PECore_DecodeAxiRead_switch_lp_mux_25_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_14_5 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl,
      rva_out_reg_data_23_17_sva_dfm_6_5, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3[5]),
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_5_0_rsp_0,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_28_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[21]),
      (rva_out_reg_data_23_17_sva_dfm_8_6_4[0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_30_nl
      = PECore_DecodeAxiRead_switch_lp_mux_28_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_14_4 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_30_nl,
      rva_out_reg_data_23_17_sva_dfm_6_4, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3[4]),
      (weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_5_0_rsp_1[4]),
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign PECore_DecodeAxiRead_switch_lp_mux_29_nl = MUX_v_4_2_2((SC_SRAM_CONFIG[20:17]),
      rva_out_reg_data_23_17_sva_dfm_8_3_0, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31_nl
      = MUX_v_4_2_2(4'b0000, PECore_DecodeAxiRead_switch_lp_mux_29_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_14_3_0 = MUX1HOT_v_4_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31_nl,
      rva_out_reg_data_23_17_sva_dfm_6_3_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3[3:0]),
      (weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_5_0_rsp_1[3:0]),
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8});
  assign weight_port_read_out_data_and_109_enex5 = weight_port_read_out_data_and_64_cse
      & reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_2_enexo;
  assign weight_port_read_out_data_and_110_enex5 = weight_port_read_out_data_and_64_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_4_2_enexo;
  assign or_dcpl_308 = weight_mem_run_3_for_5_and_159_itm_1 | weight_mem_run_3_for_5_and_158_itm_1;
  assign or_dcpl_312 = weight_mem_run_3_for_5_and_159_itm_1 | weight_mem_run_3_for_5_and_150_itm_2;
  assign or_dcpl_330 = weight_mem_run_3_for_5_and_132_itm_1 | weight_mem_run_3_for_5_and_144_itm_1;
  assign and_dcpl_719 = fsm_output & while_stage_0_7;
  assign or_dcpl_345 = weight_mem_run_3_for_5_and_94_itm_1 | weight_mem_run_3_for_5_and_92_itm_2;
  assign or_dcpl_350 = weight_mem_run_3_for_5_and_95_itm_2 | weight_mem_run_3_for_5_and_86_itm_2;
  assign or_dcpl_355 = weight_mem_run_3_for_5_and_96_itm_1 | weight_mem_run_3_for_5_and_79_itm_1;
  assign or_dcpl_382 = weight_mem_run_3_for_5_and_31_itm_2 | weight_mem_run_3_for_5_and_30_itm_2;
  assign and_dcpl_811 = while_stage_0_3 & fsm_output;
  assign or_tmp_1863 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1;
  assign data_in_tmp_operator_2_for_and_tmp = PECoreRun_wen & weight_mem_run_3_for_land_3_lpi_1_dfm_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7;
  assign pe_manager_base_input_and_tmp = PECoreRun_wen & ((or_dcpl_135 & while_stage_0_3)
      | and_dcpl_240);
  assign rva_in_reg_data_and_tmp = PECoreRun_wen & and_dcpl_297 & (and_301_cse |
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign and_2070_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b10111101) & mux_387_cse;
  assign and_2071_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b10111101);
  assign mux_742_nl = MUX_s_1_2_2(and_2070_nl, and_2071_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1656_tmp = mux_742_nl & rva_in_reg_rw_and_5_cse;
  assign and_2095_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010000))) & mux_387_cse;
  assign nor_1315_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010000));
  assign mux_780_nl = MUX_s_1_2_2(and_2095_nl, nor_1315_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1694_tmp = mux_780_nl & rva_in_reg_rw_and_5_cse;
  assign nor_801_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0001010) | mux_389_cse);
  assign nor_802_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010101));
  assign mux_406_nl = MUX_s_1_2_2(nor_801_nl, nor_802_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1320_tmp = mux_406_nl & rva_in_reg_rw_and_5_cse;
  assign and_2068_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10111100))) & mux_387_cse;
  assign nor_1261_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10111100));
  assign mux_740_nl = MUX_s_1_2_2(and_2068_nl, nor_1261_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1654_tmp = mux_740_nl & rva_in_reg_rw_and_5_cse;
  assign and_1895_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010110))) & mux_387_cse;
  assign nor_805_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010110));
  assign mux_408_nl = MUX_s_1_2_2(and_1895_nl, nor_805_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1322_tmp = mux_408_nl & rva_in_reg_rw_and_5_cse;
  assign and_2165_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11111001) & mux_387_cse;
  assign and_2166_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111001);
  assign mux_862_nl = MUX_s_1_2_2(and_2165_nl, and_2166_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1776_tmp = mux_862_nl & rva_in_reg_rw_and_5_cse;
  assign and_2113_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11011101) & mux_387_cse;
  assign and_2114_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11011101);
  assign mux_806_nl = MUX_s_1_2_2(and_2113_nl, and_2114_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1720_tmp = mux_806_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1051_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0111000) |
      mux_389_cse);
  assign nor_1052_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110001));
  assign mux_590_nl = MUX_s_1_2_2(nor_1051_nl, nor_1052_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1504_tmp = mux_590_nl & rva_in_reg_rw_and_5_cse;
  assign and_1953_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011000))) & mux_387_cse;
  assign nor_983_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011000));
  assign mux_540_nl = MUX_s_1_2_2(and_1953_nl, nor_983_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1454_tmp = mux_540_nl & rva_in_reg_rw_and_5_cse;
  assign nor_779_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0000110) | mux_389_cse);
  assign nor_780_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001101));
  assign mux_390_nl = MUX_s_1_2_2(nor_779_nl, nor_780_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1304_tmp = mux_390_nl & rva_in_reg_rw_and_5_cse;
  assign and_1900_nl = (~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[4]))
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[3])) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_818_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b000110)
      | nand_247_cse);
  assign mux_418_nl = MUX_s_1_2_2(and_1900_nl, nor_818_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1332_tmp = mux_418_nl & rva_in_reg_rw_and_5_cse;
  assign and_1939_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01001000))) & mux_387_cse;
  assign nor_941_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001000));
  assign mux_508_nl = MUX_s_1_2_2(and_1939_nl, nor_941_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1422_tmp = mux_508_nl & rva_in_reg_rw_and_5_cse;
  assign and_1914_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00101110))) & mux_387_cse;
  assign nor_869_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101110));
  assign mux_456_nl = MUX_s_1_2_2(and_1914_nl, nor_869_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1370_tmp = mux_456_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1105_nl = ~((~ (PEManager_15U_GetInputAddr_acc_tmp[7])) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[0])
      | (PEManager_15U_GetInputAddr_acc_tmp[1]) | mux_403_cse);
  assign nor_1106_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000100));
  assign mux_628_nl = MUX_s_1_2_2(nor_1105_nl, nor_1106_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1542_tmp = mux_628_nl & rva_in_reg_rw_and_5_cse;
  assign and_2028_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011011))) & mux_387_cse;
  assign nor_1167_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b100110)
      | nand_247_cse);
  assign mux_674_nl = MUX_s_1_2_2(and_2028_nl, nor_1167_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1588_tmp = mux_674_nl & rva_in_reg_rw_and_5_cse;
  assign and_2030_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011101))) & mux_387_cse;
  assign nor_1173_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011101));
  assign mux_678_nl = MUX_s_1_2_2(and_2030_nl, nor_1173_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1592_tmp = mux_678_nl & rva_in_reg_rw_and_5_cse;
  assign and_2152_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11110011) & mux_387_cse;
  assign nor_1414_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b111100)))
      | nand_247_cse);
  assign mux_850_nl = MUX_s_1_2_2(and_2152_nl, nor_1414_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1764_tmp = mux_850_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1149_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1001010) |
      mux_389_cse);
  assign nor_1150_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010101));
  assign mux_662_nl = MUX_s_1_2_2(nor_1149_nl, nor_1150_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1576_tmp = mux_662_nl & rva_in_reg_rw_and_5_cse;
  assign nor_876_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0011000) | mux_389_cse);
  assign nor_877_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110001));
  assign mux_462_nl = MUX_s_1_2_2(nor_876_nl, nor_877_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1376_tmp = mux_462_nl & rva_in_reg_rw_and_5_cse;
  assign and_2111_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11011100))) & mux_387_cse;
  assign nor_1350_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11011100));
  assign mux_804_nl = MUX_s_1_2_2(and_2111_nl, nor_1350_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1718_tmp = mux_804_nl & rva_in_reg_rw_and_5_cse;
  assign and_1954_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011010))) & mux_387_cse;
  assign nor_988_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011010));
  assign mux_544_nl = MUX_s_1_2_2(and_1954_nl, nor_988_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1458_tmp = mux_544_nl & rva_in_reg_rw_and_5_cse;
  assign and_1948_nl = (~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[6]))
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[4]))
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_969_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b010100)
      | nand_247_cse);
  assign mux_530_nl = MUX_s_1_2_2(and_1948_nl, nor_969_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1444_tmp = mux_530_nl & rva_in_reg_rw_and_5_cse;
  assign nor_963_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0101000) | mux_389_cse);
  assign nor_964_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010001));
  assign mux_526_nl = MUX_s_1_2_2(nor_963_nl, nor_964_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1440_tmp = mux_526_nl & rva_in_reg_rw_and_5_cse;
  assign and_2148_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11110001))) & mux_387_cse;
  assign nor_1408_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11110001));
  assign mux_846_nl = MUX_s_1_2_2(and_2148_nl, nor_1408_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1760_tmp = mux_846_nl & rva_in_reg_rw_and_5_cse;
  assign nor_878_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[5])) | (~ (PEManager_15U_GetInputAddr_acc_tmp[4]))
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_879_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110010));
  assign mux_464_nl = MUX_s_1_2_2(nor_878_nl, nor_879_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1378_tmp = mux_464_nl & rva_in_reg_rw_and_5_cse;
  assign and_1963_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100000))) & mux_387_cse;
  assign nor_1006_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100000));
  assign mux_556_nl = MUX_s_1_2_2(and_1963_nl, nor_1006_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1470_tmp = mux_556_nl & rva_in_reg_rw_and_5_cse;
  assign and_1995_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b01111011) & mux_387_cse;
  assign nor_1082_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b011110)))
      | nand_247_cse);
  assign mux_610_nl = MUX_s_1_2_2(and_1995_nl, nor_1082_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1524_tmp = mux_610_nl & rva_in_reg_rw_and_5_cse;
  assign and_1889_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00001100))) & mux_387_cse;
  assign nor_778_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001100));
  assign mux_388_nl = MUX_s_1_2_2(and_1889_nl, nor_778_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1302_tmp = mux_388_nl & rva_in_reg_rw_and_5_cse;
  assign and_2168_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11111010) & mux_387_cse;
  assign and_2169_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111010);
  assign mux_864_nl = MUX_s_1_2_2(and_2168_nl, and_2169_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1778_tmp = mux_864_nl & rva_in_reg_rw_and_5_cse;
  assign and_2163_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11111000))) & mux_387_cse;
  assign nor_1427_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11111000));
  assign mux_860_nl = MUX_s_1_2_2(and_2163_nl, nor_1427_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1774_tmp = mux_860_nl & rva_in_reg_rw_and_5_cse;
  assign and_2158_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11110110) & mux_387_cse;
  assign and_2159_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11110110);
  assign mux_856_nl = MUX_s_1_2_2(and_2158_nl, and_2159_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1770_tmp = mux_856_nl & rva_in_reg_rw_and_5_cse;
  assign and_1962_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b01011111) & mux_387_cse;
  assign nor_1003_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:5]!=3'b010)
      | nand_254_cse);
  assign mux_554_nl = MUX_s_1_2_2(and_1962_nl, nor_1003_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1468_tmp = mux_554_nl & rva_in_reg_rw_and_5_cse;
  assign and_2183_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11111111) & mux_387_cse;
  assign and_2184_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111111);
  assign mux_874_nl = MUX_s_1_2_2(and_2183_nl, and_2184_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1788_tmp = mux_874_nl & rva_in_reg_rw_and_5_cse;
  assign nor_791_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_792_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010001));
  assign mux_398_nl = MUX_s_1_2_2(nor_791_nl, nor_792_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1312_tmp = mux_398_nl & rva_in_reg_rw_and_5_cse;
  assign and_2136_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11101011) & mux_387_cse;
  assign nor_1392_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b111010)))
      | nand_247_cse);
  assign mux_834_nl = MUX_s_1_2_2(and_2136_nl, nor_1392_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1748_tmp = mux_834_nl & rva_in_reg_rw_and_5_cse;
  assign and_2101_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010110))) & mux_387_cse;
  assign nor_1332_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010110));
  assign mux_792_nl = MUX_s_1_2_2(and_2101_nl, nor_1332_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1706_tmp = mux_792_nl & rva_in_reg_rw_and_5_cse;
  assign and_2172_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11111011) & mux_387_cse;
  assign nor_1434_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b111110)))
      | nand_247_cse);
  assign mux_866_nl = MUX_s_1_2_2(and_2172_nl, nor_1434_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1780_tmp = mux_866_nl & rva_in_reg_rw_and_5_cse;
  assign and_2130_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11100111) & mux_387_cse;
  assign nor_1380_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b11100)
      | nand_248_cse);
  assign mux_826_nl = MUX_s_1_2_2(and_2130_nl, nor_1380_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1740_tmp = mux_826_nl & rva_in_reg_rw_and_5_cse;
  assign and_1970_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101000))) & mux_387_cse;
  assign nor_1027_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101000));
  assign mux_572_nl = MUX_s_1_2_2(and_1970_nl, nor_1027_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1486_tmp = mux_572_nl & rva_in_reg_rw_and_5_cse;
  assign and_2015_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10001110))) & mux_387_cse;
  assign nor_1132_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001110));
  assign mux_648_nl = MUX_s_1_2_2(and_2015_nl, nor_1132_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1562_tmp = mux_648_nl & rva_in_reg_rw_and_5_cse;
  assign and_1975_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101101))) & mux_387_cse;
  assign nor_1041_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101101));
  assign mux_582_nl = MUX_s_1_2_2(and_1975_nl, nor_1041_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1496_tmp = mux_582_nl & rva_in_reg_rw_and_5_cse;
  assign nor_842_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[5])) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[0])
      | (PEManager_15U_GetInputAddr_acc_tmp[1]) | mux_403_cse);
  assign nor_843_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100100));
  assign mux_436_nl = MUX_s_1_2_2(nor_842_nl, nor_843_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1350_tmp = mux_436_nl & rva_in_reg_rw_and_5_cse;
  assign or_947_nl = (state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[3]));
  assign or_945_nl = (~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[3]));
  assign mux_379_nl = MUX_s_1_2_2(or_947_nl, or_945_nl, or_898_cse);
  assign nor_765_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[2]) | (PEManager_15U_GetInputAddr_acc_tmp[0])
      | (PEManager_15U_GetInputAddr_acc_tmp[1]) | mux_379_nl);
  assign nor_766_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001000));
  assign mux_380_nl = MUX_s_1_2_2(nor_765_nl, nor_766_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1294_tmp = mux_380_nl & rva_in_reg_rw_and_5_cse;
  assign nor_797_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_798_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b000100)
      | nand_247_cse);
  assign mux_402_nl = MUX_s_1_2_2(nor_797_nl, nor_798_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1316_tmp = mux_402_nl & rva_in_reg_rw_and_5_cse;
  assign and_2057_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110101))) & mux_387_cse;
  assign nor_1240_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110101));
  assign mux_726_nl = MUX_s_1_2_2(and_2057_nl, nor_1240_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1640_tmp = mux_726_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1227_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1011000) |
      mux_389_cse);
  assign nor_1228_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110001));
  assign mux_718_nl = MUX_s_1_2_2(nor_1227_nl, nor_1228_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1632_tmp = mux_718_nl & rva_in_reg_rw_and_5_cse;
  assign and_2077_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b10111111) & mux_387_cse;
  assign nor_1268_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:6]!=2'b10)
      | nand_262_cse);
  assign mux_746_nl = MUX_s_1_2_2(and_2077_nl, nor_1268_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1660_tmp = mux_746_nl & rva_in_reg_rw_and_5_cse;
  assign nor_754_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000100) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_755_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000100));
  assign mux_372_nl = MUX_s_1_2_2(nor_754_nl, nor_755_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1286_tmp = mux_372_nl & rva_in_reg_rw_and_5_cse;
  assign and_2089_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001100))) & mux_387_cse;
  assign nor_1303_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001100));
  assign mux_772_nl = MUX_s_1_2_2(and_2089_nl, nor_1303_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1686_tmp = mux_772_nl & rva_in_reg_rw_and_5_cse;
  assign nor_886_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0011010) | mux_389_cse);
  assign nor_887_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110101));
  assign mux_470_nl = MUX_s_1_2_2(nor_886_nl, nor_887_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1384_tmp = mux_470_nl & rva_in_reg_rw_and_5_cse;
  assign and_1984_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110100))) & mux_387_cse;
  assign nor_1061_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110100));
  assign mux_596_nl = MUX_s_1_2_2(and_1984_nl, nor_1061_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1510_tmp = mux_596_nl & rva_in_reg_rw_and_5_cse;
  assign and_2013_nl = (~((~ (PEManager_15U_GetInputAddr_acc_tmp[7])) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[3])) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_1124_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b100010)
      | nand_247_cse);
  assign mux_642_nl = MUX_s_1_2_2(and_2013_nl, nor_1124_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1556_tmp = mux_642_nl & rva_in_reg_rw_and_5_cse;
  assign and_1976_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101110))) & mux_387_cse;
  assign nor_1044_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101110));
  assign mux_584_nl = MUX_s_1_2_2(and_1976_nl, nor_1044_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1498_tmp = mux_584_nl & rva_in_reg_rw_and_5_cse;
  assign and_2011_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10001000))) & mux_387_cse;
  assign nor_1117_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001000));
  assign mux_636_nl = MUX_s_1_2_2(and_2011_nl, nor_1117_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1550_tmp = mux_636_nl & rva_in_reg_rw_and_5_cse;
  assign and_1956_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011011))) & mux_387_cse;
  assign nor_991_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b010110)
      | nand_247_cse);
  assign mux_546_nl = MUX_s_1_2_2(and_1956_nl, nor_991_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1460_tmp = mux_546_nl & rva_in_reg_rw_and_5_cse;
  assign and_1923_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110111))) & mux_387_cse;
  assign nor_893_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b00110)
      | nand_248_cse);
  assign mux_474_nl = MUX_s_1_2_2(and_1923_nl, nor_893_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1388_tmp = mux_474_nl & rva_in_reg_rw_and_5_cse;
  assign nor_929_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[6]))
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[0])
      | (PEManager_15U_GetInputAddr_acc_tmp[1]) | mux_403_cse);
  assign nor_930_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000100));
  assign mux_500_nl = MUX_s_1_2_2(nor_929_nl, nor_930_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1414_tmp = mux_500_nl & rva_in_reg_rw_and_5_cse;
  assign and_2121_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100000))) & mux_387_cse;
  assign nor_1360_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100000));
  assign mux_812_nl = MUX_s_1_2_2(and_2121_nl, nor_1360_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1726_tmp = mux_812_nl & rva_in_reg_rw_and_5_cse;
  assign and_2120_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11011111) & mux_387_cse;
  assign nor_1357_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:5]==3'b110)))
      | nand_254_cse);
  assign mux_810_nl = MUX_s_1_2_2(and_2120_nl, nor_1357_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1724_tmp = mux_810_nl & rva_in_reg_rw_and_5_cse;
  assign and_1958_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011101))) & mux_387_cse;
  assign nor_997_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011101));
  assign mux_550_nl = MUX_s_1_2_2(and_1958_nl, nor_997_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1464_tmp = mux_550_nl & rva_in_reg_rw_and_5_cse;
  assign and_1941_nl = (~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[6]))
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[3])) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_948_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b010010)
      | nand_247_cse);
  assign mux_514_nl = MUX_s_1_2_2(and_1941_nl, nor_948_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1428_tmp = mux_514_nl & rva_in_reg_rw_and_5_cse;
  assign and_2010_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000111))) & mux_387_cse;
  assign nor_1114_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b10000)
      | nand_248_cse);
  assign mux_634_nl = MUX_s_1_2_2(and_2010_nl, nor_1114_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1548_tmp = mux_634_nl & rva_in_reg_rw_and_5_cse;
  assign and_2022_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010110))) & mux_387_cse;
  assign nor_1153_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010110));
  assign mux_664_nl = MUX_s_1_2_2(and_2022_nl, nor_1153_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1578_tmp = mux_664_nl & rva_in_reg_rw_and_5_cse;
  assign and_1974_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101100))) & mux_387_cse;
  assign nor_1038_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101100));
  assign mux_580_nl = MUX_s_1_2_2(and_1974_nl, nor_1038_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1494_tmp = mux_580_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1204_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1010100) |
      mux_389_cse);
  assign nor_1205_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101001));
  assign mux_702_nl = MUX_s_1_2_2(nor_1204_nl, nor_1205_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1616_tmp = mux_702_nl & rva_in_reg_rw_and_5_cse;
  assign and_1920_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110100))) & mux_387_cse;
  assign nor_885_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110100));
  assign mux_468_nl = MUX_s_1_2_2(and_1920_nl, nor_885_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1382_tmp = mux_468_nl & rva_in_reg_rw_and_5_cse;
  assign and_2147_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11110000))) & mux_387_cse;
  assign nor_1405_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11110000));
  assign mux_844_nl = MUX_s_1_2_2(and_2147_nl, nor_1405_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1758_tmp = mux_844_nl & rva_in_reg_rw_and_5_cse;
  assign and_2100_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010101))) & mux_387_cse;
  assign nor_1329_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010101));
  assign mux_790_nl = MUX_s_1_2_2(and_2100_nl, nor_1329_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1704_tmp = mux_790_nl & rva_in_reg_rw_and_5_cse;
  assign and_1991_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01111001))) & mux_387_cse;
  assign nor_1076_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111001));
  assign mux_606_nl = MUX_s_1_2_2(and_1991_nl, nor_1076_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1520_tmp = mux_606_nl & rva_in_reg_rw_and_5_cse;
  assign and_1890_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00001110))) & mux_387_cse;
  assign nor_783_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001110));
  assign mux_392_nl = MUX_s_1_2_2(and_1890_nl, nor_783_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1306_tmp = mux_392_nl & rva_in_reg_rw_and_5_cse;
  assign and_2078_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000000))) & mux_387_cse;
  assign nor_1271_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000000));
  assign mux_748_nl = MUX_s_1_2_2(and_2078_nl, nor_1271_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1662_tmp = mux_748_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1274_nl = ~((~ (PEManager_15U_GetInputAddr_acc_tmp[7])) | (~ (PEManager_15U_GetInputAddr_acc_tmp[6]))
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_1275_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000010));
  assign mux_752_nl = MUX_s_1_2_2(nor_1274_nl, nor_1275_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1666_tmp = mux_752_nl & rva_in_reg_rw_and_5_cse;
  assign and_2046_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101100))) & mux_387_cse;
  assign nor_1214_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101100));
  assign mux_708_nl = MUX_s_1_2_2(and_2046_nl, nor_1214_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1622_tmp = mux_708_nl & rva_in_reg_rw_and_5_cse;
  assign and_1985_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110101))) & mux_387_cse;
  assign nor_1064_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110101));
  assign mux_598_nl = MUX_s_1_2_2(and_1985_nl, nor_1064_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1512_tmp = mux_598_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1282_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1100010) |
      mux_389_cse);
  assign nor_1283_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000101));
  assign mux_758_nl = MUX_s_1_2_2(nor_1282_nl, nor_1283_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1672_tmp = mux_758_nl & rva_in_reg_rw_and_5_cse;
  assign and_1938_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000111))) & mux_387_cse;
  assign nor_938_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b01000)
      | nand_248_cse);
  assign mux_506_nl = MUX_s_1_2_2(and_1938_nl, nor_938_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1420_tmp = mux_506_nl & rva_in_reg_rw_and_5_cse;
  assign and_1904_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00011111))) & mux_387_cse;
  assign nor_829_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:5]!=3'b000)
      | nand_254_cse);
  assign mux_426_nl = MUX_s_1_2_2(and_1904_nl, nor_829_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1340_tmp = mux_426_nl & rva_in_reg_rw_and_5_cse;
  assign nor_855_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0010100) | mux_389_cse);
  assign nor_856_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101001));
  assign mux_446_nl = MUX_s_1_2_2(nor_855_nl, nor_856_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1360_tmp = mux_446_nl & rva_in_reg_rw_and_5_cse;
  assign and_2031_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011110))) & mux_387_cse;
  assign nor_1176_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011110));
  assign mux_680_nl = MUX_s_1_2_2(and_2031_nl, nor_1176_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1594_tmp = mux_680_nl & rva_in_reg_rw_and_5_cse;
  assign and_1925_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111010))) & mux_387_cse;
  assign nor_901_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111010));
  assign mux_480_nl = MUX_s_1_2_2(and_1925_nl, nor_901_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1394_tmp = mux_480_nl & rva_in_reg_rw_and_5_cse;
  assign and_1942_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01001100))) & mux_387_cse;
  assign nor_951_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001100));
  assign mux_516_nl = MUX_s_1_2_2(and_1942_nl, nor_951_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1430_tmp = mux_516_nl & rva_in_reg_rw_and_5_cse;
  assign and_1898_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00011000))) & mux_387_cse;
  assign nor_811_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011000));
  assign mux_412_nl = MUX_s_1_2_2(and_1898_nl, nor_811_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1326_tmp = mux_412_nl & rva_in_reg_rw_and_5_cse;
  assign nor_921_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_922_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000001));
  assign mux_494_nl = MUX_s_1_2_2(nor_921_nl, nor_922_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1408_tmp = mux_494_nl & rva_in_reg_rw_and_5_cse;
  assign and_1910_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00101000))) & mux_387_cse;
  assign nor_854_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101000));
  assign mux_444_nl = MUX_s_1_2_2(and_1910_nl, nor_854_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1358_tmp = mux_444_nl & rva_in_reg_rw_and_5_cse;
  assign and_1902_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00011110))) & mux_387_cse;
  assign nor_826_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011110));
  assign mux_424_nl = MUX_s_1_2_2(and_1902_nl, nor_826_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1338_tmp = mux_424_nl & rva_in_reg_rw_and_5_cse;
  assign and_2024_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010111))) & mux_387_cse;
  assign nor_1156_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b10010)
      | nand_248_cse);
  assign mux_666_nl = MUX_s_1_2_2(and_2024_nl, nor_1156_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1580_tmp = mux_666_nl & rva_in_reg_rw_and_5_cse;
  assign and_1913_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00101100))) & mux_387_cse;
  assign nor_864_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101100));
  assign mux_452_nl = MUX_s_1_2_2(and_1913_nl, nor_864_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1366_tmp = mux_452_nl & rva_in_reg_rw_and_5_cse;
  assign and_1973_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101011))) & mux_387_cse;
  assign nor_1035_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b011010)
      | nand_247_cse);
  assign mux_578_nl = MUX_s_1_2_2(and_1973_nl, nor_1035_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1492_tmp = mux_578_nl & rva_in_reg_rw_and_5_cse;
  assign nor_745_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_746_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000001));
  assign mux_366_nl = MUX_s_1_2_2(nor_745_nl, nor_746_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1280_tmp = mux_366_nl & rva_in_reg_rw_and_5_cse;
  assign and_1909_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100111))) & mux_387_cse;
  assign nor_851_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b00100)
      | nand_248_cse);
  assign mux_442_nl = MUX_s_1_2_2(and_1909_nl, nor_851_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1356_tmp = mux_442_nl & rva_in_reg_rw_and_5_cse;
  assign and_1929_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111101))) & mux_387_cse;
  assign nor_910_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111101));
  assign mux_486_nl = MUX_s_1_2_2(and_1929_nl, nor_910_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1400_tmp = mux_486_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1118_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1000100) |
      mux_389_cse);
  assign nor_1119_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001001));
  assign mux_638_nl = MUX_s_1_2_2(nor_1118_nl, nor_1119_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1552_tmp = mux_638_nl & rva_in_reg_rw_and_5_cse;
  assign and_2116_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11011110) & mux_387_cse;
  assign and_2117_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11011110);
  assign mux_808_nl = MUX_s_1_2_2(and_2116_nl, and_2117_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1722_tmp = mux_808_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1193_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1010010) |
      mux_389_cse);
  assign nor_1194_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100101));
  assign mux_694_nl = MUX_s_1_2_2(nor_1193_nl, nor_1194_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1608_tmp = mux_694_nl & rva_in_reg_rw_and_5_cse;
  assign and_1959_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011110))) & mux_387_cse;
  assign nor_1000_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011110));
  assign mux_552_nl = MUX_s_1_2_2(and_1959_nl, nor_1000_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1466_tmp = mux_552_nl & rva_in_reg_rw_and_5_cse;
  assign and_2180_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11111110) & mux_387_cse;
  assign and_2181_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111110);
  assign mux_872_nl = MUX_s_1_2_2(and_2180_nl, and_2181_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1786_tmp = mux_872_nl & rva_in_reg_rw_and_5_cse;
  assign and_2094_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11001111) & mux_387_cse;
  assign nor_1312_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b1100)
      | nand_250_cse);
  assign mux_778_nl = MUX_s_1_2_2(and_2094_nl, nor_1312_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1692_tmp = mux_778_nl & rva_in_reg_rw_and_5_cse;
  assign and_1916_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00101111))) & mux_387_cse;
  assign nor_872_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b0010)
      | nand_250_cse);
  assign mux_458_nl = MUX_s_1_2_2(and_1916_nl, nor_872_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1372_tmp = mux_458_nl & rva_in_reg_rw_and_5_cse;
  assign nor_984_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0101100) | mux_389_cse);
  assign nor_985_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011001));
  assign mux_542_nl = MUX_s_1_2_2(nor_984_nl, nor_985_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1456_tmp = mux_542_nl & rva_in_reg_rw_and_5_cse;
  assign and_2125_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100100))) & mux_387_cse;
  assign nor_1371_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100100));
  assign mux_820_nl = MUX_s_1_2_2(and_2125_nl, nor_1371_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1734_tmp = mux_820_nl & rva_in_reg_rw_and_5_cse;
  assign and_2133_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11101010))) & mux_387_cse;
  assign nor_1389_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11101010));
  assign mux_832_nl = MUX_s_1_2_2(and_2133_nl, nor_1389_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1746_tmp = mux_832_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1272_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1100000) |
      mux_389_cse);
  assign nor_1273_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000001));
  assign mux_750_nl = MUX_s_1_2_2(nor_1272_nl, nor_1273_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1664_tmp = mux_750_nl & rva_in_reg_rw_and_5_cse;
  assign and_2067_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b10111011) & mux_387_cse;
  assign nor_1258_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b101110)))
      | nand_247_cse);
  assign mux_738_nl = MUX_s_1_2_2(and_2067_nl, nor_1258_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1652_tmp = mux_738_nl & rva_in_reg_rw_and_5_cse;
  assign nor_865_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0010110) | mux_389_cse);
  assign nor_866_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101101));
  assign mux_454_nl = MUX_s_1_2_2(nor_865_nl, nor_866_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1368_tmp = mux_454_nl & rva_in_reg_rw_and_5_cse;
  assign and_1980_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110000))) & mux_387_cse;
  assign nor_1050_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110000));
  assign mux_588_nl = MUX_s_1_2_2(and_1980_nl, nor_1050_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1502_tmp = mux_588_nl & rva_in_reg_rw_and_5_cse;
  assign nor_774_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00001011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_775_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b000010)
      | nand_247_cse);
  assign mux_386_nl = MUX_s_1_2_2(nor_774_nl, nor_775_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1300_tmp = mux_386_nl & rva_in_reg_rw_and_5_cse;
  assign nor_924_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_925_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000010));
  assign mux_496_nl = MUX_s_1_2_2(nor_924_nl, nor_925_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1410_tmp = mux_496_nl & rva_in_reg_rw_and_5_cse;
  assign and_1892_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00001111))) & mux_387_cse;
  assign nor_786_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b0000)
      | nand_250_cse);
  assign mux_394_nl = MUX_s_1_2_2(and_1892_nl, nor_786_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1308_tmp = mux_394_nl & rva_in_reg_rw_and_5_cse;
  assign and_2062_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10111000))) & mux_387_cse;
  assign nor_1249_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10111000));
  assign mux_732_nl = MUX_s_1_2_2(and_2062_nl, nor_1249_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1646_tmp = mux_732_nl & rva_in_reg_rw_and_5_cse;
  assign and_1969_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100111))) & mux_387_cse;
  assign nor_1024_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b01100)
      | nand_248_cse);
  assign mux_570_nl = MUX_s_1_2_2(and_1969_nl, nor_1024_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1484_tmp = mux_570_nl & rva_in_reg_rw_and_5_cse;
  assign and_1996_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01111100))) & mux_387_cse;
  assign nor_1085_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111100));
  assign mux_612_nl = MUX_s_1_2_2(and_1996_nl, nor_1085_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1526_tmp = mux_612_nl & rva_in_reg_rw_and_5_cse;
  assign and_2058_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110110))) & mux_387_cse;
  assign nor_1243_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110110));
  assign mux_728_nl = MUX_s_1_2_2(and_2058_nl, nor_1243_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1642_tmp = mux_728_nl & rva_in_reg_rw_and_5_cse;
  assign and_2162_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11110111) & mux_387_cse;
  assign nor_1424_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]==5'b11110)))
      | nand_248_cse);
  assign mux_858_nl = MUX_s_1_2_2(and_2162_nl, nor_1424_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1772_tmp = mux_858_nl & rva_in_reg_rw_and_5_cse;
  assign and_1949_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010100))) & mux_387_cse;
  assign nor_972_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010100));
  assign mux_532_nl = MUX_s_1_2_2(and_1949_nl, nor_972_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1446_tmp = mux_532_nl & rva_in_reg_rw_and_5_cse;
  assign and_2041_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100111))) & mux_387_cse;
  assign nor_1200_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b10100)
      | nand_248_cse);
  assign mux_698_nl = MUX_s_1_2_2(and_2041_nl, nor_1200_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1612_tmp = mux_698_nl & rva_in_reg_rw_and_5_cse;
  assign and_2021_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010100))) & mux_387_cse;
  assign nor_1148_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010100));
  assign mux_660_nl = MUX_s_1_2_2(and_2021_nl, nor_1148_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1574_tmp = mux_660_nl & rva_in_reg_rw_and_5_cse;
  assign and_2124_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100011))) & mux_387_cse;
  assign nor_1368_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b111000)
      | nand_247_cse);
  assign mux_818_nl = MUX_s_1_2_2(and_2124_nl, nor_1368_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1732_tmp = mux_818_nl & rva_in_reg_rw_and_5_cse;
  assign and_2131_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11101000))) & mux_387_cse;
  assign nor_1383_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11101000));
  assign mux_828_nl = MUX_s_1_2_2(and_2131_nl, nor_1383_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1742_tmp = mux_828_nl & rva_in_reg_rw_and_5_cse;
  assign and_2064_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10111010))) & mux_387_cse;
  assign nor_1255_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10111010));
  assign mux_736_nl = MUX_s_1_2_2(and_2064_nl, nor_1255_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1650_tmp = mux_736_nl & rva_in_reg_rw_and_5_cse;
  assign and_2177_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11111101) & mux_387_cse;
  assign and_2178_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111101);
  assign mux_870_nl = MUX_s_1_2_2(and_2177_nl, and_2178_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1784_tmp = mux_870_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1028_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0110100) |
      mux_389_cse);
  assign nor_1029_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101001));
  assign mux_574_nl = MUX_s_1_2_2(nor_1028_nl, nor_1029_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1488_tmp = mux_574_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1017_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0110010) |
      mux_389_cse);
  assign nor_1018_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100101));
  assign mux_566_nl = MUX_s_1_2_2(nor_1017_nl, nor_1018_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1480_tmp = mux_566_nl & rva_in_reg_rw_and_5_cse;
  assign nor_763_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000111) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_764_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b00000)
      | nand_248_cse);
  assign mux_378_nl = MUX_s_1_2_2(nor_763_nl, nor_764_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1292_tmp = mux_378_nl & rva_in_reg_rw_and_5_cse;
  assign nor_757_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000101) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_758_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000101));
  assign mux_374_nl = MUX_s_1_2_2(nor_757_nl, nor_758_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1288_tmp = mux_374_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1293_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1100100) |
      mux_389_cse);
  assign nor_1294_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001001));
  assign mux_766_nl = MUX_s_1_2_2(nor_1293_nl, nor_1294_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1680_tmp = mux_766_nl & rva_in_reg_rw_and_5_cse;
  assign and_2137_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11101100))) & mux_387_cse;
  assign nor_1395_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11101100));
  assign mux_836_nl = MUX_s_1_2_2(and_2137_nl, nor_1395_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1750_tmp = mux_836_nl & rva_in_reg_rw_and_5_cse;
  assign and_2080_nl = (~((~ (PEManager_15U_GetInputAddr_acc_tmp[7])) | (~ (PEManager_15U_GetInputAddr_acc_tmp[6]))
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_1278_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b110000)
      | nand_247_cse);
  assign mux_754_nl = MUX_s_1_2_2(and_2080_nl, nor_1278_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1668_tmp = mux_754_nl & rva_in_reg_rw_and_5_cse;
  assign and_1930_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111110))) & mux_387_cse;
  assign nor_913_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111110));
  assign mux_488_nl = MUX_s_1_2_2(and_1930_nl, nor_913_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1402_tmp = mux_488_nl & rva_in_reg_rw_and_5_cse;
  assign and_1957_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011100))) & mux_387_cse;
  assign nor_994_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011100));
  assign mux_548_nl = MUX_s_1_2_2(and_1957_nl, nor_994_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1462_tmp = mux_548_nl & rva_in_reg_rw_and_5_cse;
  assign nor_794_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_795_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010010));
  assign mux_400_nl = MUX_s_1_2_2(nor_794_nl, nor_795_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1314_tmp = mux_400_nl & rva_in_reg_rw_and_5_cse;
  assign nor_840_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_841_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b001000)
      | nand_247_cse);
  assign mux_434_nl = MUX_s_1_2_2(nor_840_nl, nor_841_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1348_tmp = mux_434_nl & rva_in_reg_rw_and_5_cse;
  assign and_2096_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010010))) & mux_387_cse;
  assign nor_1320_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010010));
  assign mux_784_nl = MUX_s_1_2_2(and_2096_nl, nor_1320_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1698_tmp = mux_784_nl & rva_in_reg_rw_and_5_cse;
  assign and_1971_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101010))) & mux_387_cse;
  assign nor_1032_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101010));
  assign mux_576_nl = MUX_s_1_2_2(and_1971_nl, nor_1032_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1490_tmp = mux_576_nl & rva_in_reg_rw_and_5_cse;
  assign and_1936_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000110))) & mux_387_cse;
  assign nor_935_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000110));
  assign mux_504_nl = MUX_s_1_2_2(and_1936_nl, nor_935_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1418_tmp = mux_504_nl & rva_in_reg_rw_and_5_cse;
  assign and_2001_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b01111110) & mux_387_cse;
  assign and_2002_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b01111110);
  assign mux_616_nl = MUX_s_1_2_2(and_2001_nl, and_2002_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1530_tmp = mux_616_nl & rva_in_reg_rw_and_5_cse;
  assign input_mem_banks_read_read_data_and_30_tmp = PECoreRun_wen & and_dcpl_211;
  assign nor_751_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_752_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b000000)
      | nand_247_cse);
  assign mux_370_nl = MUX_s_1_2_2(nor_751_nl, nor_752_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1284_tmp = mux_370_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1007_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0110000) |
      mux_389_cse);
  assign nor_1008_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100001));
  assign mux_558_nl = MUX_s_1_2_2(nor_1007_nl, nor_1008_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1472_tmp = mux_558_nl & rva_in_reg_rw_and_5_cse;
  assign and_2174_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11111100) & mux_387_cse;
  assign and_2175_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111100);
  assign mux_868_nl = MUX_s_1_2_2(and_2174_nl, and_2175_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1782_tmp = mux_868_nl & rva_in_reg_rw_and_5_cse;
  assign nor_952_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0100110) | mux_389_cse);
  assign nor_953_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001101));
  assign mux_518_nl = MUX_s_1_2_2(nor_952_nl, nor_953_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1432_tmp = mux_518_nl & rva_in_reg_rw_and_5_cse;
  assign nor_897_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0011100) | mux_389_cse);
  assign nor_898_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111001));
  assign mux_478_nl = MUX_s_1_2_2(nor_897_nl, nor_898_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1392_tmp = mux_478_nl & rva_in_reg_rw_and_5_cse;
  assign and_2106_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11011001))) & mux_387_cse;
  assign nor_1341_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11011001));
  assign mux_798_nl = MUX_s_1_2_2(and_2106_nl, nor_1341_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1712_tmp = mux_798_nl & rva_in_reg_rw_and_5_cse;
  assign and_2037_nl = (~((~ (PEManager_15U_GetInputAddr_acc_tmp[7])) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[5])) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_1189_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b101000)
      | nand_247_cse);
  assign mux_690_nl = MUX_s_1_2_2(and_2037_nl, nor_1189_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1604_tmp = mux_690_nl & rva_in_reg_rw_and_5_cse;
  assign and_1893_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010000))) & mux_387_cse;
  assign nor_789_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010000));
  assign mux_396_nl = MUX_s_1_2_2(and_1893_nl, nor_789_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1310_tmp = mux_396_nl & rva_in_reg_rw_and_5_cse;
  assign nor_857_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[5])) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[3])) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_858_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101010));
  assign mux_448_nl = MUX_s_1_2_2(nor_857_nl, nor_858_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1362_tmp = mux_448_nl & rva_in_reg_rw_and_5_cse;
  assign and_2110_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11011011) & mux_387_cse;
  assign nor_1347_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b110110)))
      | nand_247_cse);
  assign mux_802_nl = MUX_s_1_2_2(and_2110_nl, nor_1347_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1716_tmp = mux_802_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1361_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1110000) |
      mux_389_cse);
  assign nor_1362_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100001));
  assign mux_814_nl = MUX_s_1_2_2(nor_1361_nl, nor_1362_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1728_tmp = mux_814_nl & rva_in_reg_rw_and_5_cse;
  assign and_1990_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01111000))) & mux_387_cse;
  assign nor_1073_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111000));
  assign mux_604_nl = MUX_s_1_2_2(and_1990_nl, nor_1073_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1518_tmp = mux_604_nl & rva_in_reg_rw_and_5_cse;
  assign and_1933_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b00111111) & mux_387_cse;
  assign nor_916_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:6]!=2'b00)
      | nand_262_cse);
  assign mux_490_nl = MUX_s_1_2_2(and_1933_nl, nor_916_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1404_tmp = mux_490_nl & rva_in_reg_rw_and_5_cse;
  assign and_2126_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100101))) & mux_387_cse;
  assign nor_1374_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100101));
  assign mux_822_nl = MUX_s_1_2_2(and_2126_nl, nor_1374_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1736_tmp = mux_822_nl & rva_in_reg_rw_and_5_cse;
  assign and_2052_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110000))) & mux_387_cse;
  assign nor_1226_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110000));
  assign mux_716_nl = MUX_s_1_2_2(and_2052_nl, nor_1226_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1630_tmp = mux_716_nl & rva_in_reg_rw_and_5_cse;
  assign and_1921_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110110))) & mux_387_cse;
  assign nor_890_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110110));
  assign mux_472_nl = MUX_s_1_2_2(and_1921_nl, nor_890_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1386_tmp = mux_472_nl & rva_in_reg_rw_and_5_cse;
  assign nor_944_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[6]))
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[3])) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_945_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001010));
  assign mux_512_nl = MUX_s_1_2_2(nor_944_nl, nor_945_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1426_tmp = mux_512_nl & rva_in_reg_rw_and_5_cse;
  assign and_1946_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010000))) & mux_387_cse;
  assign nor_962_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010000));
  assign mux_524_nl = MUX_s_1_2_2(and_1946_nl, nor_962_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1438_tmp = mux_524_nl & rva_in_reg_rw_and_5_cse;
  assign and_1943_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01001110))) & mux_387_cse;
  assign nor_956_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001110));
  assign mux_520_nl = MUX_s_1_2_2(and_1943_nl, nor_956_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1434_tmp = mux_520_nl & rva_in_reg_rw_and_5_cse;
  assign and_2014_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10001100))) & mux_387_cse;
  assign nor_1127_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001100));
  assign mux_644_nl = MUX_s_1_2_2(and_2014_nl, nor_1127_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1558_tmp = mux_644_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1160_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1001100) |
      mux_389_cse);
  assign nor_1161_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011001));
  assign mux_670_nl = MUX_s_1_2_2(nor_1160_nl, nor_1161_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1584_tmp = mux_670_nl & rva_in_reg_rw_and_5_cse;
  assign and_2048_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101110))) & mux_387_cse;
  assign nor_1220_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101110));
  assign mux_712_nl = MUX_s_1_2_2(and_2048_nl, nor_1220_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1626_tmp = mux_712_nl & rva_in_reg_rw_and_5_cse;
  assign and_2029_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011100))) & mux_387_cse;
  assign nor_1170_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011100));
  assign mux_676_nl = MUX_s_1_2_2(and_2029_nl, nor_1170_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1590_tmp = mux_676_nl & rva_in_reg_rw_and_5_cse;
  assign and_2086_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001010))) & mux_387_cse;
  assign nor_1297_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001010));
  assign mux_768_nl = MUX_s_1_2_2(and_2086_nl, nor_1297_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1682_tmp = mux_768_nl & rva_in_reg_rw_and_5_cse;
  assign and_2142_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11101110) & mux_387_cse;
  assign and_2143_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11101110);
  assign mux_840_nl = MUX_s_1_2_2(and_2142_nl, and_2143_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1754_tmp = mux_840_nl & rva_in_reg_rw_and_5_cse;
  assign nor_927_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_928_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b010000)
      | nand_247_cse);
  assign mux_498_nl = MUX_s_1_2_2(nor_927_nl, nor_928_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1412_tmp = mux_498_nl & rva_in_reg_rw_and_5_cse;
  assign and_1952_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010111))) & mux_387_cse;
  assign nor_980_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b01010)
      | nand_248_cse);
  assign mux_538_nl = MUX_s_1_2_2(and_1952_nl, nor_980_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1452_tmp = mux_538_nl & rva_in_reg_rw_and_5_cse;
  assign and_2020_nl = (~((~ (PEManager_15U_GetInputAddr_acc_tmp[7])) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[4]))
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_1145_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b100100)
      | nand_247_cse);
  assign mux_658_nl = MUX_s_1_2_2(and_2020_nl, nor_1145_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1572_tmp = mux_658_nl & rva_in_reg_rw_and_5_cse;
  assign and_2043_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101010))) & mux_387_cse;
  assign nor_1208_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101010));
  assign mux_704_nl = MUX_s_1_2_2(and_2043_nl, nor_1208_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1618_tmp = mux_704_nl & rva_in_reg_rw_and_5_cse;
  assign nor_748_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_749_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000010));
  assign mux_368_nl = MUX_s_1_2_2(nor_748_nl, nor_749_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1282_tmp = mux_368_nl & rva_in_reg_rw_and_5_cse;
  assign nor_822_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0001110) | mux_389_cse);
  assign nor_823_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011101));
  assign mux_422_nl = MUX_s_1_2_2(nor_822_nl, nor_823_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1336_tmp = mux_422_nl & rva_in_reg_rw_and_5_cse;
  assign and_2061_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b10110111) & mux_387_cse;
  assign nor_1246_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b10110)
      | nand_248_cse);
  assign mux_730_nl = MUX_s_1_2_2(and_2061_nl, nor_1246_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1644_tmp = mux_730_nl & rva_in_reg_rw_and_5_cse;
  assign and_2039_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100110))) & mux_387_cse;
  assign nor_1197_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100110));
  assign mux_696_nl = MUX_s_1_2_2(and_2039_nl, nor_1197_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1610_tmp = mux_696_nl & rva_in_reg_rw_and_5_cse;
  assign nor_834_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_835_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100001));
  assign mux_430_nl = MUX_s_1_2_2(nor_834_nl, nor_835_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1344_tmp = mux_430_nl & rva_in_reg_rw_and_5_cse;
  assign and_2008_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000110))) & mux_387_cse;
  assign nor_1111_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000110));
  assign mux_632_nl = MUX_s_1_2_2(and_2008_nl, nor_1111_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1546_tmp = mux_632_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1185_nl = ~((~ (PEManager_15U_GetInputAddr_acc_tmp[7])) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[5])) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_1186_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100010));
  assign mux_688_nl = MUX_s_1_2_2(nor_1185_nl, nor_1186_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1602_tmp = mux_688_nl & rva_in_reg_rw_and_5_cse;
  assign and_2034_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b10011111) & mux_387_cse;
  assign nor_1179_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:5]!=3'b100)
      | nand_254_cse);
  assign mux_682_nl = MUX_s_1_2_2(and_2034_nl, nor_1179_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1596_tmp = mux_682_nl & rva_in_reg_rw_and_5_cse;
  assign and_1919_nl = (~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[5])) | (~ (PEManager_15U_GetInputAddr_acc_tmp[4]))
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_882_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b001100)
      | nand_247_cse);
  assign mux_466_nl = MUX_s_1_2_2(and_1919_nl, nor_882_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1380_tmp = mux_466_nl & rva_in_reg_rw_and_5_cse;
  assign and_2025_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011000))) & mux_387_cse;
  assign nor_1159_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011000));
  assign mux_668_nl = MUX_s_1_2_2(and_2025_nl, nor_1159_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1582_tmp = mux_668_nl & rva_in_reg_rw_and_5_cse;
  assign and_2047_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101101))) & mux_387_cse;
  assign nor_1217_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101101));
  assign mux_710_nl = MUX_s_1_2_2(and_2047_nl, nor_1217_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1624_tmp = mux_710_nl & rva_in_reg_rw_and_5_cse;
  assign and_2055_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110011))) & mux_387_cse;
  assign nor_1234_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b101100)
      | nand_247_cse);
  assign mux_722_nl = MUX_s_1_2_2(and_2055_nl, nor_1234_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1636_tmp = mux_722_nl & rva_in_reg_rw_and_5_cse;
  assign and_2056_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110100))) & mux_387_cse;
  assign nor_1237_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110100));
  assign mux_724_nl = MUX_s_1_2_2(and_2056_nl, nor_1237_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1638_tmp = mux_724_nl & rva_in_reg_rw_and_5_cse;
  assign and_2018_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010000))) & mux_387_cse;
  assign nor_1138_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010000));
  assign mux_652_nl = MUX_s_1_2_2(and_2018_nl, nor_1138_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1566_tmp = mux_652_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1316_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1101000) |
      mux_389_cse);
  assign nor_1317_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010001));
  assign mux_782_nl = MUX_s_1_2_2(nor_1316_nl, nor_1317_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1696_tmp = mux_782_nl & rva_in_reg_rw_and_5_cse;
  assign and_1917_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110000))) & mux_387_cse;
  assign nor_875_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110000));
  assign mux_460_nl = MUX_s_1_2_2(and_1917_nl, nor_875_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1374_tmp = mux_460_nl & rva_in_reg_rw_and_5_cse;
  assign and_2035_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100000))) & mux_387_cse;
  assign nor_1182_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100000));
  assign mux_684_nl = MUX_s_1_2_2(and_2035_nl, nor_1182_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1598_tmp = mux_684_nl & rva_in_reg_rw_and_5_cse;
  assign and_2088_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001011))) & mux_387_cse;
  assign nor_1300_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b110010)
      | nand_247_cse);
  assign mux_770_nl = MUX_s_1_2_2(and_2088_nl, nor_1300_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1684_tmp = mux_770_nl & rva_in_reg_rw_and_5_cse;
  assign nor_799_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[4]))
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[0])
      | (PEManager_15U_GetInputAddr_acc_tmp[1]) | mux_403_cse);
  assign nor_800_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010100));
  assign mux_404_nl = MUX_s_1_2_2(nor_799_nl, nor_800_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1318_tmp = mux_404_nl & rva_in_reg_rw_and_5_cse;
  assign and_1912_nl = (~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[5])) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[3])) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_861_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b001010)
      | nand_247_cse);
  assign mux_450_nl = MUX_s_1_2_2(and_1912_nl, nor_861_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1364_tmp = mux_450_nl & rva_in_reg_rw_and_5_cse;
  assign and_2139_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11101101) & mux_387_cse;
  assign and_2140_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11101101);
  assign mux_838_nl = MUX_s_1_2_2(and_2139_nl, and_2140_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1752_tmp = mux_838_nl & rva_in_reg_rw_and_5_cse;
  assign and_1967_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100110))) & mux_387_cse;
  assign nor_1021_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100110));
  assign mux_568_nl = MUX_s_1_2_2(and_1967_nl, nor_1021_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1482_tmp = mux_568_nl & rva_in_reg_rw_and_5_cse;
  assign and_1979_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b01101111) & mux_387_cse;
  assign nor_1047_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b0110)
      | nand_250_cse);
  assign mux_586_nl = MUX_s_1_2_2(and_1979_nl, nor_1047_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1500_tmp = mux_586_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1097_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_1098_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000001));
  assign mux_622_nl = MUX_s_1_2_2(nor_1097_nl, nor_1098_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1536_tmp = mux_622_nl & rva_in_reg_rw_and_5_cse;
  assign and_1966_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100100))) & mux_387_cse;
  assign nor_1016_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100100));
  assign mux_564_nl = MUX_s_1_2_2(and_1966_nl, nor_1016_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1478_tmp = mux_564_nl & rva_in_reg_rw_and_5_cse;
  assign nor_771_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00001010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_772_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001010));
  assign mux_384_nl = MUX_s_1_2_2(nor_771_nl, nor_772_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1298_tmp = mux_384_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1139_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1001000) |
      mux_389_cse);
  assign nor_1140_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010001));
  assign mux_654_nl = MUX_s_1_2_2(nor_1139_nl, nor_1140_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1568_tmp = mux_654_nl & rva_in_reg_rw_and_5_cse;
  assign and_2146_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11101111) & mux_387_cse;
  assign nor_1402_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]==4'b1110)))
      | nand_250_cse);
  assign mux_842_nl = MUX_s_1_2_2(and_2146_nl, nor_1402_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1756_tmp = mux_842_nl & rva_in_reg_rw_and_5_cse;
  assign and_2081_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000100))) & mux_387_cse;
  assign nor_1281_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000100));
  assign mux_756_nl = MUX_s_1_2_2(and_2081_nl, nor_1281_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1670_tmp = mux_756_nl & rva_in_reg_rw_and_5_cse;
  assign and_1924_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111000))) & mux_387_cse;
  assign nor_896_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111000));
  assign mux_476_nl = MUX_s_1_2_2(and_1924_nl, nor_896_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1390_tmp = mux_476_nl & rva_in_reg_rw_and_5_cse;
  assign and_2026_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011010))) & mux_387_cse;
  assign nor_1164_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011010));
  assign mux_672_nl = MUX_s_1_2_2(and_2026_nl, nor_1164_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1586_tmp = mux_672_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1128_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1000110) |
      mux_389_cse);
  assign nor_1129_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001101));
  assign mux_646_nl = MUX_s_1_2_2(nor_1128_nl, nor_1129_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1560_tmp = mux_646_nl & rva_in_reg_rw_and_5_cse;
  assign and_2155_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11110101) & mux_387_cse;
  assign and_2156_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11110101);
  assign mux_854_nl = MUX_s_1_2_2(and_2155_nl, and_2156_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1768_tmp = mux_854_nl & rva_in_reg_rw_and_5_cse;
  assign and_2006_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000000))) & mux_387_cse;
  assign nor_1095_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000000));
  assign mux_620_nl = MUX_s_1_2_2(and_2006_nl, nor_1095_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1534_tmp = mux_620_nl & rva_in_reg_rw_and_5_cse;
  assign and_2038_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100100))) & mux_387_cse;
  assign nor_1192_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100100));
  assign mux_692_nl = MUX_s_1_2_2(and_2038_nl, nor_1192_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1606_tmp = mux_692_nl & rva_in_reg_rw_and_5_cse;
  assign and_2051_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b10101111) & mux_387_cse;
  assign nor_1223_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b1010)
      | nand_250_cse);
  assign mux_714_nl = MUX_s_1_2_2(and_2051_nl, nor_1223_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1628_tmp = mux_714_nl & rva_in_reg_rw_and_5_cse;
  assign nor_931_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0100010) | mux_389_cse);
  assign nor_932_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000101));
  assign mux_502_nl = MUX_s_1_2_2(nor_931_nl, nor_932_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1416_tmp = mux_502_nl & rva_in_reg_rw_and_5_cse;
  assign nor_760_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000110) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_761_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000110));
  assign mux_376_nl = MUX_s_1_2_2(nor_760_nl, nor_761_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1290_tmp = mux_376_nl & rva_in_reg_rw_and_5_cse;
  assign and_1998_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b01111101) & mux_387_cse;
  assign and_1999_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b01111101);
  assign mux_614_nl = MUX_s_1_2_2(and_1998_nl, and_1999_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1528_tmp = mux_614_nl & rva_in_reg_rw_and_5_cse;
  assign and_2005_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b01111111) & mux_387_cse;
  assign nor_1092_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111111));
  assign mux_618_nl = MUX_s_1_2_2(and_2005_nl, nor_1092_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1532_tmp = mux_618_nl & rva_in_reg_rw_and_5_cse;
  assign nor_965_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[6]))
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[4]))
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_966_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010010));
  assign mux_528_nl = MUX_s_1_2_2(nor_965_nl, nor_966_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1442_tmp = mux_528_nl & rva_in_reg_rw_and_5_cse;
  assign nor_812_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0001100) | mux_389_cse);
  assign nor_813_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011001));
  assign mux_414_nl = MUX_s_1_2_2(nor_812_nl, nor_813_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1328_tmp = mux_414_nl & rva_in_reg_rw_and_5_cse;
  assign and_2122_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100010))) & mux_387_cse;
  assign nor_1365_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100010));
  assign mux_816_nl = MUX_s_1_2_2(and_2122_nl, nor_1365_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1730_tmp = mux_816_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1120_nl = ~((~ (PEManager_15U_GetInputAddr_acc_tmp[7])) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[3])) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_1121_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001010));
  assign mux_640_nl = MUX_s_1_2_2(nor_1120_nl, nor_1121_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1554_tmp = mux_640_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1107_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1000010) |
      mux_389_cse);
  assign nor_1108_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000101));
  assign mux_630_nl = MUX_s_1_2_2(nor_1107_nl, nor_1108_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1544_tmp = mux_630_nl & rva_in_reg_rw_and_5_cse;
  assign nor_844_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0010010) | mux_389_cse);
  assign nor_845_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100101));
  assign mux_438_nl = MUX_s_1_2_2(nor_844_nl, nor_845_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1352_tmp = mux_438_nl & rva_in_reg_rw_and_5_cse;
  assign and_2149_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11110010))) & mux_387_cse;
  assign nor_1411_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11110010));
  assign mux_848_nl = MUX_s_1_2_2(and_2149_nl, nor_1411_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1762_tmp = mux_848_nl & rva_in_reg_rw_and_5_cse;
  assign and_2045_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101011))) & mux_387_cse;
  assign nor_1211_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b101010)
      | nand_247_cse);
  assign mux_706_nl = MUX_s_1_2_2(and_2045_nl, nor_1211_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1620_tmp = mux_706_nl & rva_in_reg_rw_and_5_cse;
  assign and_2105_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11011000))) & mux_387_cse;
  assign nor_1338_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11011000));
  assign mux_796_nl = MUX_s_1_2_2(and_2105_nl, nor_1338_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1710_tmp = mux_796_nl & rva_in_reg_rw_and_5_cse;
  assign and_2091_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001110))) & mux_387_cse;
  assign nor_1309_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001110));
  assign mux_776_nl = MUX_s_1_2_2(and_2091_nl, nor_1309_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1690_tmp = mux_776_nl & rva_in_reg_rw_and_5_cse;
  assign nor_768_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00001001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_769_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001001));
  assign mux_382_nl = MUX_s_1_2_2(nor_768_nl, nor_769_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1296_tmp = mux_382_nl & rva_in_reg_rw_and_5_cse;
  assign and_1905_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100000))) & mux_387_cse;
  assign nor_832_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100000));
  assign mux_428_nl = MUX_s_1_2_2(and_1905_nl, nor_832_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1342_tmp = mux_428_nl & rva_in_reg_rw_and_5_cse;
  assign and_1950_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010110))) & mux_387_cse;
  assign nor_977_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010110));
  assign mux_536_nl = MUX_s_1_2_2(and_1950_nl, nor_977_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1450_tmp = mux_536_nl & rva_in_reg_rw_and_5_cse;
  assign and_1992_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01111010))) & mux_387_cse;
  assign nor_1079_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111010));
  assign mux_608_nl = MUX_s_1_2_2(and_1992_nl, nor_1079_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1522_tmp = mux_608_nl & rva_in_reg_rw_and_5_cse;
  assign nor_814_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[4]))
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[3])) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_815_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011010));
  assign mux_416_nl = MUX_s_1_2_2(nor_814_nl, nor_815_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1330_tmp = mux_416_nl & rva_in_reg_rw_and_5_cse;
  assign and_2073_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b10111110) & mux_387_cse;
  assign and_2074_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b10111110);
  assign mux_744_nl = MUX_s_1_2_2(and_2073_nl, and_2074_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1658_tmp = mux_744_nl & rva_in_reg_rw_and_5_cse;
  assign and_2084_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000111))) & mux_387_cse;
  assign nor_1289_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b11000)
      | nand_248_cse);
  assign mux_762_nl = MUX_s_1_2_2(and_2084_nl, nor_1289_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1676_tmp = mux_762_nl & rva_in_reg_rw_and_5_cse;
  assign nor_942_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0100100) | mux_389_cse);
  assign nor_943_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001001));
  assign mux_510_nl = MUX_s_1_2_2(nor_942_nl, nor_943_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1424_tmp = mux_510_nl & rva_in_reg_rw_and_5_cse;
  assign and_1945_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01001111))) & mux_387_cse;
  assign nor_959_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b0100)
      | nand_250_cse);
  assign mux_522_nl = MUX_s_1_2_2(and_1945_nl, nor_959_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1436_tmp = mux_522_nl & rva_in_reg_rw_and_5_cse;
  assign and_1981_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110010))) & mux_387_cse;
  assign nor_1055_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110010));
  assign mux_592_nl = MUX_s_1_2_2(and_1981_nl, nor_1055_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1506_tmp = mux_592_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1103_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_1104_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b100000)
      | nand_247_cse);
  assign mux_626_nl = MUX_s_1_2_2(nor_1103_nl, nor_1104_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1540_tmp = mux_626_nl & rva_in_reg_rw_and_5_cse;
  assign and_2082_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000110))) & mux_387_cse;
  assign nor_1286_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000110));
  assign mux_760_nl = MUX_s_1_2_2(and_2082_nl, nor_1286_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1674_tmp = mux_760_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1009_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[6]))
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[5])) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_1010_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100010));
  assign mux_560_nl = MUX_s_1_2_2(nor_1009_nl, nor_1010_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1474_tmp = mux_560_nl & rva_in_reg_rw_and_5_cse;
  assign and_2042_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101000))) & mux_387_cse;
  assign nor_1203_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101000));
  assign mux_700_nl = MUX_s_1_2_2(and_2042_nl, nor_1203_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1614_tmp = mux_700_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1141_nl = ~((~ (PEManager_15U_GetInputAddr_acc_tmp[7])) | (PEManager_15U_GetInputAddr_acc_tmp[6])
      | (PEManager_15U_GetInputAddr_acc_tmp[5]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[4]))
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (PEManager_15U_GetInputAddr_acc_tmp[0]) | mux_415_cse);
  assign nor_1142_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010010));
  assign mux_656_nl = MUX_s_1_2_2(nor_1141_nl, nor_1142_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1570_tmp = mux_656_nl & rva_in_reg_rw_and_5_cse;
  assign and_2098_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010011))) & mux_387_cse;
  assign nor_1323_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b110100)
      | nand_247_cse);
  assign mux_786_nl = MUX_s_1_2_2(and_2098_nl, nor_1323_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1700_tmp = mux_786_nl & rva_in_reg_rw_and_5_cse;
  assign and_2132_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11101001))) & mux_387_cse;
  assign nor_1386_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11101001));
  assign mux_830_nl = MUX_s_1_2_2(and_2132_nl, nor_1386_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1744_tmp = mux_830_nl & rva_in_reg_rw_and_5_cse;
  assign and_1983_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110011))) & mux_387_cse;
  assign nor_1058_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b011100)
      | nand_247_cse);
  assign mux_594_nl = MUX_s_1_2_2(and_1983_nl, nor_1058_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1508_tmp = mux_594_nl & rva_in_reg_rw_and_5_cse;
  assign and_2104_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11010111) & mux_387_cse;
  assign nor_1335_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b11010)
      | nand_248_cse);
  assign mux_794_nl = MUX_s_1_2_2(and_2104_nl, nor_1335_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1708_tmp = mux_794_nl & rva_in_reg_rw_and_5_cse;
  assign and_2099_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010100))) & mux_387_cse;
  assign nor_1326_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010100));
  assign mux_788_nl = MUX_s_1_2_2(and_2099_nl, nor_1326_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1702_tmp = mux_788_nl & rva_in_reg_rw_and_5_cse;
  assign and_2085_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001000))) & mux_387_cse;
  assign nor_1292_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001000));
  assign mux_764_nl = MUX_s_1_2_2(and_2085_nl, nor_1292_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1678_tmp = mux_764_nl & rva_in_reg_rw_and_5_cse;
  assign and_2017_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10001111))) & mux_387_cse;
  assign nor_1135_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b1000)
      | nand_250_cse);
  assign mux_650_nl = MUX_s_1_2_2(and_2017_nl, nor_1135_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1564_tmp = mux_650_nl & rva_in_reg_rw_and_5_cse;
  assign and_2063_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10111001))) & mux_387_cse;
  assign nor_1252_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10111001));
  assign mux_734_nl = MUX_s_1_2_2(and_2063_nl, nor_1252_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1648_tmp = mux_734_nl & rva_in_reg_rw_and_5_cse;
  assign and_1897_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010111))) & mux_387_cse;
  assign nor_808_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b00010)
      | nand_248_cse);
  assign mux_410_nl = MUX_s_1_2_2(and_1897_nl, nor_808_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1324_tmp = mux_410_nl & rva_in_reg_rw_and_5_cse;
  assign and_2090_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001101))) & mux_387_cse;
  assign nor_1306_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001101));
  assign mux_774_nl = MUX_s_1_2_2(and_2090_nl, nor_1306_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1688_tmp = mux_774_nl & rva_in_reg_rw_and_5_cse;
  assign and_1965_nl = (~((PEManager_15U_GetInputAddr_acc_tmp[7]) | (~ (PEManager_15U_GetInputAddr_acc_tmp[6]))
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[5])) | (PEManager_15U_GetInputAddr_acc_tmp[4])
      | (PEManager_15U_GetInputAddr_acc_tmp[3]) | (PEManager_15U_GetInputAddr_acc_tmp[2])
      | (~ (PEManager_15U_GetInputAddr_acc_tmp[0])))) & mux_417_cse;
  assign nor_1013_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b011000)
      | nand_247_cse);
  assign mux_562_nl = MUX_s_1_2_2(and_1965_nl, nor_1013_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1476_tmp = mux_562_nl & rva_in_reg_rw_and_5_cse;
  assign and_1907_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100110))) & mux_387_cse;
  assign nor_848_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100110));
  assign mux_440_nl = MUX_s_1_2_2(and_1907_nl, nor_848_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1354_tmp = mux_440_nl & rva_in_reg_rw_and_5_cse;
  assign and_2127_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100110))) & mux_387_cse;
  assign nor_1377_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100110));
  assign mux_824_nl = MUX_s_1_2_2(and_2127_nl, nor_1377_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1738_tmp = mux_824_nl & rva_in_reg_rw_and_5_cse;
  assign and_2107_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11011010))) & mux_387_cse;
  assign nor_1344_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11011010));
  assign mux_800_nl = MUX_s_1_2_2(and_2107_nl, nor_1344_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1714_tmp = mux_800_nl & rva_in_reg_rw_and_5_cse;
  assign and_2153_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11110100))) & mux_387_cse;
  assign nor_1417_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11110100));
  assign mux_852_nl = MUX_s_1_2_2(and_2153_nl, nor_1417_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1766_tmp = mux_852_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1183_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1010000) |
      mux_389_cse);
  assign nor_1184_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100001));
  assign mux_686_nl = MUX_s_1_2_2(nor_1183_nl, nor_1184_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1600_tmp = mux_686_nl & rva_in_reg_rw_and_5_cse;
  assign and_1928_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111100))) & mux_387_cse;
  assign nor_907_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111100));
  assign mux_484_nl = MUX_s_1_2_2(and_1928_nl, nor_907_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1398_tmp = mux_484_nl & rva_in_reg_rw_and_5_cse;
  assign nor_1100_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_1101_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000010));
  assign mux_624_nl = MUX_s_1_2_2(nor_1100_nl, nor_1101_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1538_tmp = mux_624_nl & rva_in_reg_rw_and_5_cse;
  assign and_2053_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110010))) & mux_387_cse;
  assign nor_1231_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110010));
  assign mux_720_nl = MUX_s_1_2_2(and_2053_nl, nor_1231_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1634_tmp = mux_720_nl & rva_in_reg_rw_and_5_cse;
  assign and_1989_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b01110111) & mux_387_cse;
  assign nor_1070_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b01110)
      | nand_248_cse);
  assign mux_602_nl = MUX_s_1_2_2(and_1989_nl, nor_1070_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1516_tmp = mux_602_nl & rva_in_reg_rw_and_5_cse;
  assign and_1986_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110110))) & mux_387_cse;
  assign nor_1067_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110110));
  assign mux_600_nl = MUX_s_1_2_2(and_1986_nl, nor_1067_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1514_tmp = mux_600_nl & rva_in_reg_rw_and_5_cse;
  assign nor_837_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_365_cse));
  assign nor_838_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100010));
  assign mux_432_nl = MUX_s_1_2_2(nor_837_nl, nor_838_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1346_tmp = mux_432_nl & rva_in_reg_rw_and_5_cse;
  assign and_1901_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00011100))) & mux_387_cse;
  assign nor_821_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011100));
  assign mux_420_nl = MUX_s_1_2_2(and_1901_nl, nor_821_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1334_tmp = mux_420_nl & rva_in_reg_rw_and_5_cse;
  assign nor_973_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0101010) | mux_389_cse);
  assign nor_974_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010101));
  assign mux_534_nl = MUX_s_1_2_2(nor_973_nl, nor_974_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1448_tmp = mux_534_nl & rva_in_reg_rw_and_5_cse;
  assign and_1934_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000000))) & mux_387_cse;
  assign nor_919_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000000));
  assign mux_492_nl = MUX_s_1_2_2(and_1934_nl, nor_919_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1406_tmp = mux_492_nl & rva_in_reg_rw_and_5_cse;
  assign and_1927_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111011))) & mux_387_cse;
  assign nor_904_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b001110)
      | nand_247_cse);
  assign mux_482_nl = MUX_s_1_2_2(and_1927_nl, nor_904_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1396_tmp = mux_482_nl & rva_in_reg_rw_and_5_cse;
  assign or_900_nl = (state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1;
  assign or_899_nl = (~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1;
  assign mux_363_nl = MUX_s_1_2_2(or_900_nl, or_899_nl, or_898_cse);
  assign nor_742_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000000) | mux_363_nl);
  assign nor_743_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000000));
  assign mux_364_nl = MUX_s_1_2_2(nor_742_nl, nor_743_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1278_tmp = mux_364_nl & rva_in_reg_rw_and_5_cse;
  assign input_mem_banks_read_read_data_and_29_tmp = PECoreRun_wen & (~((~((~ rva_in_reg_rw_sva_st_1_4)
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)))
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
      & while_stage_0_6;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_31_cse <= 1'b0;
      reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_21_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_act_port_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      pe_config_manager_counter_sva_dfm_3_1 <= 4'b0000;
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= 1'b0;
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= 1'b0;
      while_stage_0_3 <= 1'b0;
      while_stage_0_4 <= 1'b0;
      while_stage_0_5 <= 1'b0;
      while_stage_0_6 <= 1'b0;
      while_stage_0_7 <= 1'b0;
      while_stage_0_8 <= 1'b0;
      while_stage_0_9 <= 1'b0;
      while_stage_0_10 <= 1'b0;
      while_stage_0_11 <= 1'b0;
      while_stage_0_12 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_1_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1
          <= 1'b0;
      input_read_addrs_sva_1_1 <= 8'b00000000;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= 1'b0;
    end
    else if ( PECoreRun_wen ) begin
      reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_31_cse <= and_489_rmff;
      reg_Datapath_for_4_ProductSum_for_acc_5_cmp_cgo_ir_21_cse <= and_492_rmff;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= and_497_rmff;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= and_502_rmff;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= and_505_rmff;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= and_508_rmff;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= and_511_rmff;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= and_514_rmff;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= and_517_rmff;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= and_520_rmff;
      reg_rva_out_Push_mioi_iswt0_cse <= and_522_cse;
      reg_start_PopNB_mioi_iswt0_cse <= and_524_rmff;
      reg_act_port_Push_mioi_iswt0_cse <= and_526_rmff;
      reg_rva_in_PopNB_mioi_iswt0_cse <= fsm_output;
      pe_config_manager_counter_sva_dfm_3_1 <= MUX_v_4_2_2(4'b0000, operator_4_false_acc_nl,
          pe_config_UpdateManagerCounter_if_not_7_nl);
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= ~((pe_config_input_counter_sva_mx1 != (operator_16_false_acc_sdt_sva_1[7:0]))
          | (operator_16_false_acc_sdt_sva_1[8]));
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
      while_stage_0_3 <= reg_rva_in_PopNB_mioi_iswt0_cse;
      while_stage_0_4 <= while_stage_0_3;
      while_stage_0_5 <= while_stage_0_4;
      while_stage_0_6 <= while_stage_0_5;
      while_stage_0_7 <= while_stage_0_6;
      while_stage_0_8 <= while_stage_0_7;
      while_stage_0_9 <= while_stage_0_8;
      while_stage_0_10 <= while_stage_0_9;
      while_stage_0_11 <= while_stage_0_10;
      while_stage_0_12 <= while_stage_0_11;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[1];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1 <= pe_manager_base_weight_sva_mx2[2];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[0];
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_1_itm_1 <= ~ (pe_manager_base_weight_sva_mx1_3_0[1]);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= (pe_manager_base_weight_sva_mx2[2])
          & (pe_manager_base_weight_sva_mx1_3_0[1:0]==2'b01) & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1
          <= ~((pe_manager_base_weight_sva_mx2[2]) | (pe_manager_base_weight_sva_mx1_3_0[1:0]!=2'b00));
      input_read_addrs_sva_1_1 <= nl_input_read_addrs_sva_1_1[7:0];
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_10 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_2_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_10 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_10 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_10 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_8 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_90_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_8 <= rva_out_reg_data_30_25_sva_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_63_sva_dfm_4_5 <= 1'b0;
      rva_out_reg_data_47_sva_dfm_4_5 <= 1'b0;
      input_read_req_valid_lpi_1_dfm_1_10 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8 <= 1'b0;
      rva_out_reg_data_46_40_sva_dfm_4_5_6_4 <= 3'b000;
      rva_out_reg_data_39_36_sva_dfm_4_5_3 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_5_2 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_5_1_0 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_17_cse ) begin
      rva_out_reg_data_63_sva_dfm_4_5 <= rva_out_reg_data_63_sva_dfm_4_4;
      rva_out_reg_data_47_sva_dfm_4_5 <= rva_out_reg_data_47_sva_dfm_4_4;
      input_read_req_valid_lpi_1_dfm_1_10 <= input_read_req_valid_lpi_1_dfm_1_9;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
      rva_out_reg_data_46_40_sva_dfm_4_5_6_4 <= reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd;
      rva_out_reg_data_39_36_sva_dfm_4_5_3 <= reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd;
      rva_out_reg_data_39_36_sva_dfm_4_5_2 <= reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1;
      rva_out_reg_data_39_36_sva_dfm_4_5_1_0 <= reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_91_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_5 <= rva_out_reg_data_62_56_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_5 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_92_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_5 <= rva_out_reg_data_35_32_sva_dfm_4_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_3 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_6 <=
          1'b0;
      weight_port_read_out_data_0_3_sva_dfm_5_7 <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_6 <=
          1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_6 <=
          1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_5_0_rsp_0
          <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_5_6_0_rsp_0 <= 3'b000;
    end
    else if ( weight_port_read_out_data_and_64_cse ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2 <= weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2 <= weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2 <= weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_6 <=
          reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd;
      weight_port_read_out_data_0_3_sva_dfm_5_7 <= reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_6 <=
          reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_6 <=
          reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_5_0_rsp_0
          <= reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_1_ftd;
      weight_port_read_out_data_0_3_sva_dfm_5_6_0_rsp_0 <= reg_weight_port_read_out_data_0_3_sva_dfm_4_1_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_7_1_sva_dfm_6_6 <= 1'b0;
      rva_out_reg_data_7_1_sva_dfm_6_5_0 <= 6'b000000;
      rva_out_reg_data_15_9_sva_dfm_6_6 <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_6_5_0 <= 6'b000000;
      rva_out_reg_data_30_25_sva_dfm_6_5_3 <= 3'b000;
      rva_out_reg_data_30_25_sva_dfm_6_2_0 <= 3'b000;
      rva_out_reg_data_0_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_8_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_16_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_31_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_24_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_6_6 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_6_5 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_6_4 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_6_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_cse ) begin
      rva_out_reg_data_7_1_sva_dfm_6_6 <= PECore_PushAxiRsp_if_mux1h_10_6;
      rva_out_reg_data_7_1_sva_dfm_6_5_0 <= PECore_PushAxiRsp_if_mux1h_10_5_0;
      rva_out_reg_data_15_9_sva_dfm_6_6 <= PECore_PushAxiRsp_if_mux1h_12_6;
      rva_out_reg_data_15_9_sva_dfm_6_5_0 <= PECore_PushAxiRsp_if_mux1h_12_5_0;
      rva_out_reg_data_30_25_sva_dfm_6_5_3 <= PECore_PushAxiRsp_if_mux1h_16_5_3;
      rva_out_reg_data_30_25_sva_dfm_6_2_0 <= PECore_PushAxiRsp_if_mux1h_16_2_0;
      rva_out_reg_data_0_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_14_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
      rva_out_reg_data_8_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_15_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
      rva_out_reg_data_16_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_16_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_2, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_8);
      rva_out_reg_data_31_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_17;
      rva_out_reg_data_24_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_15;
      rva_out_reg_data_23_17_sva_dfm_6_6 <= PECore_PushAxiRsp_if_mux1h_14_6;
      rva_out_reg_data_23_17_sva_dfm_6_5 <= PECore_PushAxiRsp_if_mux1h_14_5;
      rva_out_reg_data_23_17_sva_dfm_6_4 <= PECore_PushAxiRsp_if_mux1h_14_4;
      rva_out_reg_data_23_17_sva_dfm_6_3_0 <= PECore_PushAxiRsp_if_mux1h_14_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_31_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_32_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_33_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_34_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_3
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_10 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
          <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_cse ) begin
      rva_in_reg_rw_sva_10 <= rva_in_reg_rw_sva_9;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_10 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_4 ) begin
      rva_in_reg_rw_sva_st_1_10 <= rva_in_reg_rw_sva_st_1_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_10
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_10
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_15_0_sva_dfm_1_2 <= 16'b0000000000000000;
    end
    else if ( act_port_reg_data_and_30_enex5 ) begin
      act_port_reg_data_15_0_sva_dfm_1_2 <= act_port_reg_data_15_0_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_239_224_sva_dfm_1_2 <= 16'b0000000000000000;
    end
    else if ( act_port_reg_data_and_31_enex5 ) begin
      act_port_reg_data_239_224_sva_dfm_1_2 <= act_port_reg_data_239_224_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_47_32_sva_dfm_1_2 <= 16'b0000000000000000;
    end
    else if ( act_port_reg_data_and_32_enex5 ) begin
      act_port_reg_data_47_32_sva_dfm_1_2 <= act_port_reg_data_47_32_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_207_192_sva_dfm_1_2 <= 16'b0000000000000000;
    end
    else if ( act_port_reg_data_and_33_enex5 ) begin
      act_port_reg_data_207_192_sva_dfm_1_2 <= act_port_reg_data_207_192_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_79_64_sva_dfm_1_1 <= 16'b0000000000000000;
    end
    else if ( (PECore_UpdateFSM_switch_lp_equal_tmp_2_10 | (~ while_stage_0_12) |
        while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10
        | (PECore_RunScale_PECore_RunScale_if_and_1_svs_9 & (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_9)))
        & rva_in_reg_rw_and_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)
        & ((~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9) | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9)
        ) begin
      act_port_reg_data_79_64_sva_dfm_1_1 <= MUX_v_16_2_2((readslicef_27_16_11(PECore_RunScale_if_for_3_scaled_val_mul_1_nl)),
          act_port_reg_data_79_64_sva_mx1, or_418_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_175_160_sva_dfm_1_2 <= 16'b0000000000000000;
    end
    else if ( act_port_reg_data_and_34_enex5 ) begin
      act_port_reg_data_175_160_sva_dfm_1_2 <= act_port_reg_data_175_160_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_111_96_sva_dfm_1_2 <= 16'b0000000000000000;
    end
    else if ( act_port_reg_data_and_35_enex5 ) begin
      act_port_reg_data_111_96_sva_dfm_1_2 <= act_port_reg_data_111_96_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_143_128_sva_dfm_1_2 <= 16'b0000000000000000;
    end
    else if ( act_port_reg_data_and_36_enex5 ) begin
      act_port_reg_data_143_128_sva_dfm_1_2 <= act_port_reg_data_143_128_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_10 <= 1'b0;
    end
    else if ( PECore_PushOutput_if_and_cse ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_10 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_10 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_9 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_9 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_9 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= 1'b0;
      rva_in_reg_rw_sva_9 <= 1'b0;
    end
    else if ( while_if_and_6_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
      rva_in_reg_rw_sva_9 <= rva_in_reg_rw_sva_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_8 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_27 ) begin
      rva_in_reg_rw_sva_st_1_8 <= rva_in_reg_rw_sva_st_1_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_1_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_8 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= 1'b0;
      rva_in_reg_rw_sva_8 <= 1'b0;
    end
    else if ( while_if_and_7_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
      rva_in_reg_rw_sva_8 <= rva_in_reg_rw_sva_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_30 ) begin
      rva_in_reg_rw_sva_st_1_7 <= rva_in_reg_rw_sva_st_1_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_2_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= 1'b0;
      rva_in_reg_rw_sva_7 <= 1'b0;
    end
    else if ( while_if_and_8_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
      rva_in_reg_rw_sva_7 <= rva_in_reg_rw_sva_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_enex5 ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= 1'b0;
      rva_in_reg_rw_sva_6 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_cse ) begin
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= weight_mem_run_3_for_land_3_lpi_1_dfm_2;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
      rva_in_reg_rw_sva_6 <= rva_in_reg_rw_sva_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_3_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_5,
          weight_port_read_out_data_0_7_sva_dfm_3_7, PECore_PushAxiRsp_if_else_mux_13_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_24_cse , while_and_23_cse});
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5,
          (weight_port_read_out_data_0_5_sva_dfm_3_7_4[3]), PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_24_cse , while_and_23_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & while_stage_0_6 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & while_stage_0_6 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_5 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_43 ) begin
      rva_in_reg_rw_sva_st_1_5 <= rva_in_reg_rw_sva_st_1_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1 <= 1'b0;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_156_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_158_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_159_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_144_itm_1 <= 1'b0;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_run_3_for_5_and_103_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2 <= 1'b0;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_92_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_94_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_95_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_96_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_84_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_86_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_79_itm_1 <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_28_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_30_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_31_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_20_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_22_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_23_itm_1 <= 1'b0;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= 1'b0;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_run_3_for_5_and_8_itm_1 <= 1'b0;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_162_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_163_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_164_itm_2 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_165_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_166_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_167_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_168_itm_2_cse <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= 1'b0;
    end
    else if ( weight_mem_banks_read_1_read_data_and_8_cse ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= MUX_v_64_2_2(weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= MUX_v_64_2_2(weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= MUX_v_64_2_2(weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_19_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_2_2_0!=3'b000));
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_156_itm_2 <= weight_mem_run_3_for_5_and_156_itm_1;
      weight_mem_run_3_for_5_and_158_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_159_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_150_itm_2 <= weight_mem_run_3_for_5_and_150_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1;
      weight_mem_run_3_for_5_and_144_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b111)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= weight_read_addrs_7_lpi_1_dfm_2_2_0;
      weight_mem_run_3_for_5_and_103_itm_2 <= weight_mem_run_3_for_5_and_103_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_1;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_92_itm_2 <= weight_mem_run_3_for_5_and_92_itm_1;
      weight_mem_run_3_for_5_and_94_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b101)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_95_itm_2 <= weight_mem_run_3_for_5_and_95_itm_1;
      weight_mem_run_3_for_5_and_96_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b111)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1 <= ~((weight_read_addrs_5_lpi_1_dfm_2_2_0!=3'b000));
      weight_mem_run_3_for_5_and_84_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b011)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_86_itm_2 <= weight_mem_run_3_for_5_and_86_itm_1;
      weight_mem_run_3_for_5_and_79_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b110)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= weight_read_addrs_5_lpi_1_dfm_2_2_0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1_1;
      weight_mem_run_3_for_5_and_28_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1_1;
      weight_mem_run_3_for_5_and_30_itm_2 <= weight_mem_run_3_for_5_and_30_itm_1;
      weight_mem_run_3_for_5_and_31_itm_2 <= weight_mem_run_3_for_5_and_31_itm_1;
      weight_mem_run_3_for_5_and_20_itm_2 <= weight_mem_run_3_for_5_and_20_itm_1;
      weight_mem_run_3_for_5_and_22_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1;
      weight_mem_run_3_for_5_and_23_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= weight_read_addrs_3_lpi_1_dfm_2_2_0;
      weight_mem_run_3_for_5_and_8_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1;
      reg_weight_mem_run_3_for_5_and_162_itm_2_cse <= weight_mem_run_3_for_5_and_162_itm_1;
      reg_weight_mem_run_3_for_5_and_163_itm_2_cse <= weight_mem_run_3_for_5_and_163_itm_1;
      weight_mem_run_3_for_5_and_164_itm_2 <= weight_mem_run_3_for_5_and_164_itm_1;
      reg_weight_mem_run_3_for_5_and_165_itm_2_cse <= weight_mem_run_3_for_5_and_165_itm_1;
      reg_weight_mem_run_3_for_5_and_166_itm_2_cse <= weight_mem_run_3_for_5_and_166_itm_1;
      reg_weight_mem_run_3_for_5_and_167_itm_2_cse <= weight_mem_run_3_for_5_and_167_itm_1;
      reg_weight_mem_run_3_for_5_and_168_itm_2_cse <= weight_mem_run_3_for_5_and_168_itm_1;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & while_stage_0_6 & weight_mem_run_3_for_land_3_lpi_1_dfm_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_6_nl & while_stage_0_6 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= 1'b0;
    end
    else if ( PECoreRun_wen & while_stage_0_6 & weight_mem_run_3_for_land_5_lpi_1_dfm_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2 <= 2'b00;
    end
    else if ( PECoreRun_wen & mux_8_nl & while_stage_0_6 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_2 <= MUX_v_2_2_2(pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_2[7:6]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & weight_mem_run_3_for_land_7_lpi_1_dfm_1 & while_stage_0_6
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_9_nl & while_stage_0_6 ) begin
      reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_8_itm_2_cse <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_2_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_132_itm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= 1'b0;
      rva_in_reg_rw_sva_5 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_1_cse ) begin
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= weight_mem_run_3_for_land_1_lpi_1_dfm_2;
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= weight_mem_run_3_for_land_7_lpi_1_dfm_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= weight_mem_run_3_for_land_3_lpi_1_dfm_1;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= weight_mem_run_3_for_land_5_lpi_1_dfm_1;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_132_itm_1 <= MUX_s_1_2_2(weight_mem_run_3_for_5_and_100_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
      rva_in_reg_rw_sva_5 <= rva_in_reg_rw_sva_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_71_cse ) begin
      weight_port_read_out_data_6_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_7_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_10_cse ) begin
      weight_port_read_out_data_1_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
      weight_port_read_out_data_1_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
      weight_port_read_out_data_1_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
      weight_port_read_out_data_1_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
      weight_port_read_out_data_1_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005;
      weight_port_read_out_data_1_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004;
      weight_port_read_out_data_1_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006;
      weight_port_read_out_data_1_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_000000;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_18_cse ) begin
      weight_port_read_out_data_2_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
      weight_port_read_out_data_2_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
      weight_port_read_out_data_2_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004;
      weight_port_read_out_data_2_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
      weight_port_read_out_data_2_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005;
      weight_port_read_out_data_2_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_sva_1;
      weight_port_read_out_data_2_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_6_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_7_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_24_cse ) begin
      weight_port_read_out_data_4_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_3_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_32_cse ) begin
      weight_port_read_out_data_3_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
      weight_port_read_out_data_3_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
      weight_port_read_out_data_3_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
      weight_port_read_out_data_3_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_7_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1010_cse | or_dcpl_308 | weight_mem_run_3_for_5_and_156_itm_2)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_7_sva_dfm_1 <= weight_port_read_out_data_7_7_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1010_cse | or_dcpl_312 | weight_mem_run_3_for_5_and_156_itm_2)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_6_sva_dfm_1 <= weight_port_read_out_data_7_6_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_3_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1019_cse ) begin
      weight_port_read_out_data_7_5_sva_dfm_1 <= weight_port_read_out_data_7_5_sva_dfm_2;
      weight_port_read_out_data_7_3_sva_dfm_1 <= weight_port_read_out_data_7_3_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_4_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1010_cse | or_dcpl_312 | weight_mem_run_3_for_5_and_132_itm_1)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_4_sva_dfm_1 <= weight_port_read_out_data_7_4_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_2_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1030_cse | or_dcpl_312 | or_dcpl_330) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_2_sva_dfm_1 <= weight_port_read_out_data_7_2_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1018_cse | or_dcpl_308 | or_dcpl_330) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_1_sva_dfm_1 <= weight_port_read_out_data_7_1_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1030_cse | weight_mem_run_3_for_5_and_144_itm_1 | weight_mem_run_3_for_5_and_103_itm_2
        | weight_mem_run_3_for_5_and_150_itm_2 | weight_mem_run_3_for_5_and_132_itm_1)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_0_sva_dfm_1 <= weight_port_read_out_data_7_0_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1044_cse ) begin
      weight_port_read_out_data_5_7_sva_dfm_1 <= weight_port_read_out_data_5_7_sva_dfm_3;
      weight_port_read_out_data_5_0_sva_dfm_1 <= weight_port_read_out_data_5_0_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (((xor_7_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1)
        & weight_mem_run_3_for_land_6_lpi_1_dfm_2) | or_dcpl_350 | weight_mem_run_3_for_5_and_84_itm_1)
        & and_dcpl_719 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_5_6_sva_dfm_1 <= weight_port_read_out_data_5_6_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_3_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1054_cse ) begin
      weight_port_read_out_data_5_5_sva_dfm_1 <= weight_port_read_out_data_5_5_sva_dfm_3;
      weight_port_read_out_data_5_3_sva_dfm_1 <= weight_port_read_out_data_5_3_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_2_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1059_cse ) begin
      weight_port_read_out_data_5_4_sva_dfm_1 <= weight_port_read_out_data_5_4_sva_dfm_3;
      weight_port_read_out_data_5_2_sva_dfm_1 <= weight_port_read_out_data_5_2_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1043_cse | or_dcpl_355 | weight_mem_run_3_for_5_and_86_itm_2 |
        weight_mem_run_3_for_5_and_92_itm_2) & and_dcpl_719 & PECoreRun_wen & (~
        while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_5_1_sva_dfm_1 <= weight_port_read_out_data_5_1_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_7_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1083_cse | or_dcpl_382 | weight_mem_run_3_for_5_and_28_itm_1)
        & and_dcpl_719 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_3_7_sva_dfm_1 <= weight_port_read_out_data_3_7_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1083_cse | weight_mem_run_3_for_5_and_23_itm_1 | weight_mem_run_3_for_5_and_22_itm_1
        | weight_mem_run_3_for_5_and_20_itm_2) & and_dcpl_719 & PECoreRun_wen & (~
        while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_3_6_sva_dfm_1 <= weight_port_read_out_data_3_6_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_5_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (((xor_13_cse | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse)
        & weight_mem_run_3_for_land_4_lpi_1_dfm_2) | or_dcpl_382 | weight_mem_run_3_for_5_and_20_itm_2)
        & and_dcpl_719 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_3_5_sva_dfm_1 <= weight_port_read_out_data_3_5_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_4_sva_dfm_1 <= 8'b00000000;
    end
    else if ( ((((((weight_read_addrs_3_lpi_1_dfm_3_2_0[2:1]!=2'b00)) ^ (weight_read_addrs_3_lpi_1_dfm_3_2_0[0]))
        | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse) & weight_mem_run_3_for_land_4_lpi_1_dfm_2)
        | weight_mem_run_3_for_5_and_8_itm_1 | weight_mem_run_3_for_5_and_30_itm_2
        | weight_mem_run_3_for_5_and_20_itm_2) & and_dcpl_719 & PECoreRun_wen & (~
        while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      weight_port_read_out_data_3_4_sva_dfm_1 <= weight_port_read_out_data_3_4_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_31_nl & while_stage_0_6 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_101_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 <= 1'b0;
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_113_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_itm_mx0w1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_20_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_116_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= 8'b00000000;
    end
    else if ( (weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_32_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= MUX_v_8_2_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[7:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_33_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= MUX_v_8_2_2((weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[7:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_63_8 <= 56'b00000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_218 | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & mux_35_nl ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_63_8 <= weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63:8];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_218 | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & mux_37_nl ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_RunFSM_switch_lp_equal_tmp_1_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_UpdateFSM_switch_lp_equal_tmp_2_3 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_empty_sva_1[2])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_38_nl) & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_7_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_882_cse & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_74 & and_882_cse ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= 1'b0;
      rva_in_reg_rw_sva_4 <= 1'b0;
    end
    else if ( while_if_and_11_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_87_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 | and_713_cse
          | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp
          | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp
          | and_715_cse | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp
          | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & or_296_cse;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= weight_mem_run_3_for_weight_mem_run_3_for_and_4_cse;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & or_286_cse;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
      rva_in_reg_rw_sva_4 <= rva_in_reg_rw_sva_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_49_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_55_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_61_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= weight_mem_read_arbxbar_arbiters_next_5_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_67_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_73_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_79_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_85_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse & (and_882_cse | Arbiter_8U_Roundrobin_pick_and_12_cse)
        & or_dcpl_68 ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0,
          Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1, Arbiter_8U_Roundrobin_pick_and_12_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_91_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva <= 15'b000000000000000;
    end
    else if ( (~ mux_360_nl) & fsm_output & while_stage_0_5 & PECoreRun_wen ) begin
      pe_manager_base_weight_sva <= pe_manager_base_weight_sva_mx2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= 11'b00000000000;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= 1'b0;
    end
    else if ( weight_read_addrs_and_9_cse ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= MUX_v_11_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl,
          weight_read_addrs_0_14_4_lpi_1_dfm_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= MUX_s_1_2_2((weight_read_addrs_0_3_0_lpi_1_dfm_4[3]),
          (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_24_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_25_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_26_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_27_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_28_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_29_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_30_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_31_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= 12'b000000000000;
    end
    else if ( weight_write_addrs_and_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= weight_write_addrs_lpi_1_dfm_1_2[14:3];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_153 & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]))
        ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= 1'b0;
      weight_read_addrs_1_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_3_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= 13'b0000000000000;
      weight_read_addrs_5_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_7_lpi_1_dfm_1 <= 15'b000000000000000;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1,
          and_142_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1,
          and_142_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1,
          and_142_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1,
          and_142_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1,
          and_142_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1,
          and_142_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1,
          and_142_cse);
      weight_read_addrs_1_lpi_1_dfm_1 <= weight_read_addrs_1_lpi_1_dfm_1_1;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_3_lpi_1_dfm_1 <= weight_read_addrs_3_lpi_1_dfm_1_1;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_1 <= weight_read_addrs_5_lpi_1_dfm_1_1;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_7_lpi_1_dfm_1 <= weight_read_addrs_7_lpi_1_dfm_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_23_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_1_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
          & Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_1_tmp;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_not_185,
          weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0, and_dcpl_544);
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0, and_107_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0, and_114_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0, and_121_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0, and_128_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0, and_135_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0,
          (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_1_tmp);
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0, and_142_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= 1'b0;
      rva_in_reg_rw_sva_3 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= 1'b0;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      rva_in_reg_rw_sva_3 <= reg_rva_in_reg_rw_sva_2_cse;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_23_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= 8'b00000000;
      rva_in_reg_rw_sva_st_1_3 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_55_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= 1'b0;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= 8'b00000000;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_1_for_and_cse ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
      rva_in_reg_rw_sva_st_1_3 <= reg_rva_in_reg_rw_sva_2_cse;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_55_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b101)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b011)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b110)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= weight_mem_write_arbxbar_xbar_for_lshift_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_and_75_cse ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_545);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_545);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_545);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_545);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_545);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_545);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_545);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_545);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_64_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse & ((~ while_stage_0_5) | while_and_1126_itm_1)
        ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= MUX_v_15_2_2(pe_manager_base_weight_sva_mx2,
          PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1, while_and_1126_itm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_32_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_7_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_33_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_6_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_34_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_5_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_35_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_36_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_3_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_37_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_2_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_38_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_1_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_39_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= 15'b000000000000000;
    end
    else if ( weight_write_addrs_and_2_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= pe_manager_base_input_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( weight_write_data_data_and_8_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_2_cse <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= 1'b0;
      while_and_1126_itm_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_5_cse ) begin
      reg_rva_in_reg_rw_sva_2_cse <= reg_rva_in_reg_rw_sva_st_1_1_cse;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= MUX_s_1_2_2(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
      while_and_1126_itm_1 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1
          & PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
          & reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= 4'b0000;
    end
    else if ( weight_read_addrs_and_28_enex5 ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= 11'b00000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_198 ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_2_1_sva <= 2'b00;
      pe_config_is_zero_first_sva <= 1'b0;
    end
    else if ( state_and_cse ) begin
      state_2_1_sva <= state_mux_1_cse;
      pe_config_is_zero_first_sva <= pe_config_is_zero_first_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_0_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_228) ) begin
      state_0_sva <= PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_manager_counter_sva <= 4'b0000;
    end
    else if ( (((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4:2]!=3'b000))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:5]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10:8]!=3'b000))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:11]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
        & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])
        & rva_in_PopNB_mioi_return_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]==2'b00)
        & and_dcpl_203) | and_1109_cse) & PECoreRun_wen ) begin
      pe_config_manager_counter_sva <= MUX_v_4_2_2(pe_config_manager_counter_sva_dfm_3_1,
          PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl,
          and_600_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_num_manager_sva <= 4'b0001;
      pe_config_num_output_sva <= 8'b00000001;
    end
    else if ( pe_config_num_manager_and_cse ) begin
      pe_config_num_manager_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[35:32];
      pe_config_num_output_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= 1'b0;
      state_2_1_sva_dfm_1 <= 2'b00;
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= 8'b00000000;
      input_write_req_valid_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_6_cse ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= rva_in_PopNB_mioi_return_rsc_z_mxwt;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
      state_2_1_sva_dfm_1 <= MUX_v_2_2_2(PECore_UpdateFSM_switch_lp_and_1_nl, state_mux_1_cse,
          rva_in_PopNB_mioi_return_rsc_z_mxwt);
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= and_301_cse;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0];
      input_write_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= 1'b0;
      PECore_RunFSM_switch_lp_nor_tmp_1 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_9_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= PECore_UpdateFSM_switch_lp_equal_tmp_6;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= ~(PECore_RunScale_PECore_RunScale_if_and_1_svs_1
          | PECore_UpdateFSM_switch_lp_nor_tmp_1);
      PECore_RunFSM_switch_lp_nor_tmp_1 <= ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
          | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(or_220_cse | or_dcpl_228 | (~ fsm_output))) & (mux_142_cse
        | rva_in_PopNB_mioi_return_rsc_z_mxwt | (~ reg_rva_in_PopNB_mioi_iswt0_cse))
        ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= input_port_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva <= 8'b00000000;
    end
    else if ( or_835_cse & mux_361_nl & and_dcpl_811 & PECoreRun_wen ) begin
      pe_config_input_counter_sva <= pe_config_input_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva <= 8'b00000000;
    end
    else if ( or_835_cse & mux_362_nl & and_dcpl_811 & PECoreRun_wen ) begin
      pe_config_output_counter_sva <= pe_config_output_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      operator_8_false_acc_sdt_sva_1 <= 9'b000000000;
    end
    else if ( pe_config_UpdateManagerCounter_if_if_and_enex5 ) begin
      operator_8_false_acc_sdt_sva_1 <= nl_operator_8_false_acc_sdt_sva_1[8:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiWrite_switch_lp_and_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_79_64_sva <= 16'b0000000000000000;
    end
    else if ( or_228_cse_1 & fsm_output & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_10)
        & while_stage_0_12 ) begin
      act_port_reg_data_79_64_sva <= act_port_reg_data_79_64_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_2_18_0_sva <= 19'b0000000000000000000;
    end
    else if ( (PECore_RunMac_PECore_RunMac_if_and_svs_st_9 | PECore_UpdateFSM_switch_lp_equal_tmp_2_9)
        & while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)
        & PECoreRun_wen ) begin
      accum_vector_data_2_18_0_sva <= MUX_v_19_2_2(19'b0000000000000000000, ProductSum_for_acc_21_nl,
          PECore_UpdateFSM_switch_lp_not_19_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_129_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_115_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_122_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_94_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_108_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_6_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_130_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_131_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_133_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~ mux_tmp_60) & and_dcpl_43 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
        ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= MUX_v_8_2_2(8'b00000000, mux1h_1_nl, not_2217_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_9_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_123_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_126_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[23:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_127_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[15:8]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_128_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_10_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_109_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_110_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_112_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[15:8]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_114_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~ mux_68_nl) & while_stage_0_6 ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= MUX_v_8_2_2(8'b00000000, mux_321_nl, nor_425_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_14_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_124_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_125_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_16_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_132_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[7:0]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_78_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_19_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_111_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[23:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_113_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= 1'b0;
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_5_and_156_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_150_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_103_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_95_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_92_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_86_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_31_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_30_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_20_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_168_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_167_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_166_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_165_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_164_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_163_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_162_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= 1'b0;
    end
    else if ( weight_read_addrs_and_19_cse ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= weight_read_addrs_7_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= weight_read_addrs_5_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= weight_read_addrs_3_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_5_and_156_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_150_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_17_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_103_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_95_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b110)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_92_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_11_itm_1 <= ~((weight_read_addrs_5_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_86_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b101)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_31_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1_1;
      weight_mem_run_3_for_5_and_30_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1;
      weight_mem_run_3_for_5_and_20_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= ~((weight_read_addrs_3_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_168_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
      weight_mem_run_3_for_5_and_167_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
      weight_mem_run_3_for_5_and_166_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b101)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_165_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
      weight_mem_run_3_for_5_and_164_itm_1 <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          & (pe_manager_base_weight_sva[0]) & (~ (pe_manager_base_weight_sva[2]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_163_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
      weight_mem_run_3_for_5_and_162_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1 <= ~((pe_manager_base_weight_sva[2:0]!=3'b000));
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_71_nl ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        | (~ while_stage_0_6))) ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~((~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        | (~ while_stage_0_6))) ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_73_nl ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_74_nl ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & mux_75_nl ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_24_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_29_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= 1'b0;
    end
    else if ( operator_15_false_1_and_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_142_cse | or_dcpl_59)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_or_1_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        | (~ while_stage_0_4))) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_135_cse | or_dcpl_59)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_128_cse | or_dcpl_59)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_121_cse | or_dcpl_59)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_114_cse | or_dcpl_59)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_107_cse | or_dcpl_59)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= 15'b000000000000000;
    end
    else if ( PEManager_15U_PEManagerWrite_and_enex5 ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= rva_in_reg_data_sva_1[30:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_num_input_sva <= 8'b00000001;
      pe_manager_base_bias_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_num_input_and_cse ) begin
      pe_manager_num_input_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      pe_manager_base_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[46:32];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_is_valid_sva <= 1'b0;
      pe_config_is_cluster_sva <= 1'b0;
      pe_config_is_bias_sva <= 1'b0;
    end
    else if ( pe_config_is_valid_and_cse ) begin
      pe_config_is_valid_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
      pe_config_is_cluster_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[16];
      pe_config_is_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_zero_active_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & and_301_cse & (~ PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)
        & (~ or_dcpl_239) ) begin
      pe_manager_zero_active_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva_dfm_1 <= 8'b00000000;
      pe_config_input_counter_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1169_cse ) begin
      pe_config_output_counter_sva_dfm_1 <= MUX_v_8_2_2(8'b00000000, pe_config_output_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
      pe_config_input_counter_sva_dfm_1 <= MUX_v_8_2_2(8'b00000000, pe_config_input_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_mux_19_itm_1 <= 1'b0;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= 4'b0000;
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= 11'b00000000000;
    end
    else if ( while_if_and_15_cse ) begin
      while_if_mux_19_itm_1 <= MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_19_nl,
          rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:0])
          & ({{3{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_4_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:4])
          & ({{10{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_11_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_4 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_7_cse ) begin
      rva_in_reg_rw_sva_st_1_4 <= rva_in_reg_rw_sva_st_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & PECore_PushAxiRsp_and_2_cse ) begin
      rva_in_reg_rw_sva_st_1_6 <= rva_in_reg_rw_sva_st_1_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_9 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_244 ) begin
      rva_in_reg_rw_sva_st_1_9 <= rva_in_reg_rw_sva_st_1_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= 4'b0000;
      input_read_req_valid_lpi_1_dfm_1_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= 1'b0;
    end
    else if ( while_if_and_16_cse ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16];
      input_read_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= (pe_config_num_output_sva[7]) & (~(and_301_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1))
          & PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_1 <= 2'b00;
    end
    else if ( PECoreRun_wen & or_261_cse & and_dcpl_248 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_7_itm_1 <= pe_manager_base_weight_sva[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_122_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_55_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_128_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_24_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= MUX_v_3_2_2((weight_read_addrs_1_lpi_1_dfm_1[2:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse
        & and_dcpl_248 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1
          <= ~((weight_read_addrs_1_lpi_1_dfm_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2
          <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_74_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b011)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1 <= (pe_manager_base_weight_sva[2])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1 & (pe_manager_base_weight_sva[0])
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1
          & (pe_manager_base_weight_sva[1:0]==2'b10) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1 <= (pe_manager_base_weight_sva[2])
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 & (~ (pe_manager_base_weight_sva[1]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1
          & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 & (~ (pe_manager_base_weight_sva[1]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1
          <= ~(pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1 | (pe_manager_base_weight_sva[1:0]!=2'b00));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_79_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_25_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[7]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_nl,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_23_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[5]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_22_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[4]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_1[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          PECore_UpdateFSM_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_nl,
          PECore_RunFSM_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_76_nl & while_stage_0_5 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          input_read_req_valid_lpi_1_dfm_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1 <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd
          <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1 <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd
          <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1 <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd
          <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_1_ftd
          <= 1'b0;
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd <= 1'b0;
      reg_weight_port_read_out_data_0_3_sva_dfm_4_1_ftd <= 3'b000;
    end
    else if ( weight_port_read_out_data_and_79_cse ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1 <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1[0];
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd
          <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1 <= weight_port_read_out_data_0_1_sva_dfm_3_rsp_1[0];
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd
          <= weight_port_read_out_data_0_1_sva_dfm_3_rsp_0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1 <= weight_port_read_out_data_0_2_sva_dfm_3_rsp_1_rsp_1[0];
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd
          <= weight_port_read_out_data_0_2_sva_dfm_3_rsp_0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_1_ftd
          <= weight_port_read_out_data_0_2_sva_dfm_3_rsp_1_rsp_0;
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd <= weight_port_read_out_data_0_3_sva_dfm_3_rsp_0;
      reg_weight_port_read_out_data_0_3_sva_dfm_4_1_ftd <= weight_port_read_out_data_0_3_sva_dfm_3_rsp_1_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_9_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1
          <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_95_enex5 ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1
          <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1[6:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_35_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1
          <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_96_enex5 ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1
          <= weight_port_read_out_data_0_1_sva_dfm_3_rsp_1[6:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_36_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_1_ftd_1
          <= 5'b00000;
    end
    else if ( weight_port_read_out_data_and_97_enex5 ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_1_ftd_1
          <= weight_port_read_out_data_0_2_sva_dfm_3_rsp_1_rsp_1[5:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_37_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_38_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_15_0_sva_dfm_1_1 <= 16'b0000000000000000;
      act_port_reg_data_47_32_sva_dfm_1_1 <= 16'b0000000000000000;
      act_port_reg_data_111_96_sva_dfm_1_1 <= 16'b0000000000000000;
      act_port_reg_data_143_128_sva_dfm_1_1 <= 16'b0000000000000000;
      act_port_reg_data_175_160_sva_dfm_1_1 <= 16'b0000000000000000;
      act_port_reg_data_207_192_sva_dfm_1_1 <= 16'b0000000000000000;
      act_port_reg_data_239_224_sva_dfm_1_1 <= 16'b0000000000000000;
    end
    else if ( and_1197_cse ) begin
      act_port_reg_data_15_0_sva_dfm_1_1 <= MUX_v_16_2_2((readslicef_27_16_11(PECore_RunScale_if_for_1_scaled_val_mul_1_nl)),
          act_port_reg_data_15_0_sva_mx1, or_dcpl_278);
      act_port_reg_data_47_32_sva_dfm_1_1 <= MUX_v_16_2_2((readslicef_27_16_11(PECore_RunScale_if_for_2_scaled_val_mul_1_nl)),
          act_port_reg_data_47_32_sva_mx1, or_dcpl_278);
      act_port_reg_data_111_96_sva_dfm_1_1 <= MUX_v_16_2_2((readslicef_27_16_11(PECore_RunScale_if_for_4_scaled_val_mul_1_nl)),
          act_port_reg_data_111_96_sva_mx1, or_dcpl_278);
      act_port_reg_data_143_128_sva_dfm_1_1 <= MUX_v_16_2_2((readslicef_27_16_11(PECore_RunScale_if_for_5_scaled_val_mul_1_nl)),
          act_port_reg_data_143_128_sva_mx1, or_dcpl_278);
      act_port_reg_data_175_160_sva_dfm_1_1 <= MUX_v_16_2_2((readslicef_27_16_11(PECore_RunScale_if_for_6_scaled_val_mul_1_nl)),
          act_port_reg_data_175_160_sva_mx1, or_dcpl_278);
      act_port_reg_data_207_192_sva_dfm_1_1 <= MUX_v_16_2_2((readslicef_27_16_11(PECore_RunScale_if_for_7_scaled_val_mul_1_nl)),
          act_port_reg_data_207_192_sva_mx1, or_dcpl_278);
      act_port_reg_data_239_224_sva_dfm_1_1 <= MUX_v_16_2_2((readslicef_27_16_11(PECore_RunScale_if_for_8_scaled_val_mul_1_nl)),
          act_port_reg_data_239_224_sva_mx1, or_dcpl_278);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & or_286_cse & and_dcpl_248 ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_78_nl) & while_stage_0_5 ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= MUX_s_1_2_2((weight_read_addrs_4_14_2_lpi_1_dfm_1[0]),
          weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & or_296_cse & and_dcpl_248 ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_9 <= 1'b0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd <= 1'b0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1 <= 1'b0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_2 <= 2'b00;
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd <= 3'b000;
      rva_out_reg_data_47_sva_dfm_4_4 <= 1'b0;
      rva_out_reg_data_63_sva_dfm_4_4 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( input_read_req_valid_and_1_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_9 <= input_read_req_valid_lpi_1_dfm_1_8;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd <= rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_2 <= rva_out_reg_data_39_36_sva_dfm_4_3_rsp_2;
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd <= rva_out_reg_data_46_40_sva_dfm_4_3_rsp_0;
      rva_out_reg_data_47_sva_dfm_4_4 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      rva_out_reg_data_63_sva_dfm_4_4 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_8;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_7_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_93_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= rva_out_reg_data_30_25_sva_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_ftd <= 3'b000;
      reg_rva_out_reg_data_15_9_sva_dfm_9_ftd <= 1'b0;
    end
    else if ( rva_out_reg_data_and_24_cse ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_ftd <= rva_out_reg_data_23_17_sva_dfm_6_rsp_0;
      reg_rva_out_reg_data_15_9_sva_dfm_9_ftd <= rva_out_reg_data_15_9_sva_dfm_8_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_ftd_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_94_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_ftd_1 <= rva_out_reg_data_23_17_sva_dfm_6_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_ftd_1 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_95_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_ftd_1 <= rva_out_reg_data_15_9_sva_dfm_8_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_1_ftd_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_98_enex5 ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_1_ftd_1 <= weight_port_read_out_data_0_3_sva_dfm_3_rsp_1_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_96_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= rva_out_reg_data_35_32_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_97_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_46_40_sva_dfm_4_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_98_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_4 <= rva_out_reg_data_62_56_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_99_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd <= rva_out_reg_data_55_48_sva_dfm_4_3_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_100_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_55_48_sva_dfm_4_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_15_0_sva <= 16'b0000000000000000;
      act_port_reg_data_47_32_sva <= 16'b0000000000000000;
      act_port_reg_data_111_96_sva <= 16'b0000000000000000;
      act_port_reg_data_143_128_sva <= 16'b0000000000000000;
      act_port_reg_data_175_160_sva <= 16'b0000000000000000;
      act_port_reg_data_207_192_sva <= 16'b0000000000000000;
      act_port_reg_data_239_224_sva <= 16'b0000000000000000;
    end
    else if ( and_1231_cse ) begin
      act_port_reg_data_15_0_sva <= act_port_reg_data_15_0_sva_mx1;
      act_port_reg_data_47_32_sva <= act_port_reg_data_47_32_sva_mx1;
      act_port_reg_data_111_96_sva <= act_port_reg_data_111_96_sva_mx1;
      act_port_reg_data_143_128_sva <= act_port_reg_data_143_128_sva_mx1;
      act_port_reg_data_175_160_sva <= act_port_reg_data_175_160_sva_mx1;
      act_port_reg_data_207_192_sva <= act_port_reg_data_207_192_sva_mx1;
      act_port_reg_data_239_224_sva <= act_port_reg_data_239_224_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_acc_22_itm_1 <= 19'b0000000000000000000;
      Datapath_for_3_ProductSum_for_acc_3_1 <= 18'b000000000000000000;
    end
    else if ( ProductSum_for_and_cse ) begin
      ProductSum_for_acc_22_itm_1 <= nl_ProductSum_for_acc_22_itm_1[18:0];
      Datapath_for_3_ProductSum_for_acc_3_1 <= Datapath_for_4_ProductSum_for_acc_5_cmp_22_z;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_18_0_sva <= 19'b0000000000000000000;
      accum_vector_data_0_18_0_sva <= 19'b0000000000000000000;
      accum_vector_data_6_18_0_sva <= 19'b0000000000000000000;
      accum_vector_data_1_18_0_sva <= 19'b0000000000000000000;
      accum_vector_data_5_18_0_sva <= 19'b0000000000000000000;
      accum_vector_data_4_18_0_sva <= 19'b0000000000000000000;
      accum_vector_data_3_18_0_sva <= 19'b0000000000000000000;
    end
    else if ( and_1258_cse ) begin
      accum_vector_data_7_18_0_sva <= MUX_v_19_2_2(19'b0000000000000000000, ProductSum_for_acc_nl,
          PECore_UpdateFSM_switch_lp_not_32_nl);
      accum_vector_data_0_18_0_sva <= MUX_v_19_2_2(19'b0000000000000000000, ProductSum_for_acc_33_nl,
          PECore_UpdateFSM_switch_lp_not_21_nl);
      accum_vector_data_6_18_0_sva <= MUX_v_19_2_2(19'b0000000000000000000, ProductSum_for_acc_30_nl,
          PECore_UpdateFSM_switch_lp_not_33_nl);
      accum_vector_data_1_18_0_sva <= MUX_v_19_2_2(19'b0000000000000000000, ProductSum_for_acc_27_nl,
          PECore_UpdateFSM_switch_lp_not_37_nl);
      accum_vector_data_5_18_0_sva <= MUX_v_19_2_2(19'b0000000000000000000, ProductSum_for_acc_24_nl,
          PECore_UpdateFSM_switch_lp_not_34_nl);
      accum_vector_data_4_18_0_sva <= MUX_v_19_2_2(19'b0000000000000000000, ProductSum_for_acc_18_nl,
          PECore_UpdateFSM_switch_lp_not_35_nl);
      accum_vector_data_3_18_0_sva <= MUX_v_19_2_2(19'b0000000000000000000, ProductSum_for_acc_15_nl,
          PECore_UpdateFSM_switch_lp_not_36_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_1_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= 8'b00000000;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_empty_and_enex5 ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= weight_mem_write_arbxbar_xbar_for_empty_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_data_sva_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rva_in_reg_data_and_tmp ) begin
      rva_in_reg_data_sva_1 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_18_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[0];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[8];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[16];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[31];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_39_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[7:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_40_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[15:9];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_41_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[23:17];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_42_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[30:25];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_2 <= 2'b00;
      rva_out_reg_data_46_40_sva_dfm_4_3_rsp_0 <= 3'b000;
    end
    else if ( input_read_req_valid_and_2_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= input_read_req_valid_lpi_1_dfm_1_7;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_39_36_sva_dfm_4_2_3;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_39_36_sva_dfm_4_2_2;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_2 <= rva_out_reg_data_39_36_sva_dfm_4_2_1_0;
      rva_out_reg_data_46_40_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_46_40_sva_dfm_4_2_6_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_11_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_6 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_101_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_6 <= rva_out_reg_data_30_25_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_102_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= rva_out_reg_data_35_32_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_103_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_3 <= rva_out_reg_data_62_56_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_27_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0 <= input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_6_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= MUX_v_64_2_2(input_mem_banks_read_1_for_mux_4_nl,
          input_mem_banks_read_read_data_sva_1, and_633_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_2_3 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_2_2 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_2_1_0 <= 2'b00;
      rva_out_reg_data_46_40_sva_dfm_4_2_6_4 <= 3'b000;
    end
    else if ( input_read_req_valid_and_3_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= input_read_req_valid_lpi_1_dfm_1_6;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
      rva_out_reg_data_39_36_sva_dfm_4_2_3 <= rva_out_reg_data_39_36_sva_dfm_4_1_3;
      rva_out_reg_data_39_36_sva_dfm_4_2_2 <= rva_out_reg_data_39_36_sva_dfm_4_1_2;
      rva_out_reg_data_39_36_sva_dfm_4_2_1_0 <= rva_out_reg_data_39_36_sva_dfm_4_1_1_0;
      rva_out_reg_data_46_40_sva_dfm_4_2_6_4 <= rva_out_reg_data_46_40_sva_dfm_4_1_6_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_15_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_104_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= rva_out_reg_data_30_25_sva_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_105_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= rva_out_reg_data_35_32_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_106_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_2 <= rva_out_reg_data_62_56_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_2_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1278_tmp ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= input_mem_banks_bank_a_0_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1280_tmp ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= input_mem_banks_bank_a_1_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1282_tmp ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= input_mem_banks_bank_a_2_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1284_tmp ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= input_mem_banks_bank_a_3_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1286_tmp ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= input_mem_banks_bank_a_4_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1288_tmp ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= input_mem_banks_bank_a_5_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1290_tmp ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= input_mem_banks_bank_a_6_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1292_tmp ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= input_mem_banks_bank_a_7_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1294_tmp ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= input_mem_banks_bank_a_8_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1296_tmp ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= input_mem_banks_bank_a_9_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1298_tmp ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= input_mem_banks_bank_a_10_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1300_tmp ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= input_mem_banks_bank_a_11_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1302_tmp ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= input_mem_banks_bank_a_12_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1304_tmp ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= input_mem_banks_bank_a_13_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1306_tmp ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= input_mem_banks_bank_a_14_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1308_tmp ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= input_mem_banks_bank_a_15_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1310_tmp ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= input_mem_banks_bank_a_16_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1312_tmp ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= input_mem_banks_bank_a_17_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1314_tmp ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= input_mem_banks_bank_a_18_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1316_tmp ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= input_mem_banks_bank_a_19_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1318_tmp ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= input_mem_banks_bank_a_20_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1320_tmp ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= input_mem_banks_bank_a_21_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1322_tmp ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= input_mem_banks_bank_a_22_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1324_tmp ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= input_mem_banks_bank_a_23_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1326_tmp ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= input_mem_banks_bank_a_24_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1328_tmp ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= input_mem_banks_bank_a_25_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1330_tmp ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= input_mem_banks_bank_a_26_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1332_tmp ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= input_mem_banks_bank_a_27_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1334_tmp ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= input_mem_banks_bank_a_28_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1336_tmp ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= input_mem_banks_bank_a_29_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1338_tmp ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= input_mem_banks_bank_a_30_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1340_tmp ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= input_mem_banks_bank_a_31_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1342_tmp ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= input_mem_banks_bank_a_32_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1344_tmp ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= input_mem_banks_bank_a_33_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1346_tmp ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= input_mem_banks_bank_a_34_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1348_tmp ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= input_mem_banks_bank_a_35_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1350_tmp ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= input_mem_banks_bank_a_36_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1352_tmp ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= input_mem_banks_bank_a_37_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1354_tmp ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= input_mem_banks_bank_a_38_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1356_tmp ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= input_mem_banks_bank_a_39_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1358_tmp ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= input_mem_banks_bank_a_40_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1360_tmp ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= input_mem_banks_bank_a_41_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1362_tmp ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= input_mem_banks_bank_a_42_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1364_tmp ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= input_mem_banks_bank_a_43_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1366_tmp ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= input_mem_banks_bank_a_44_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1368_tmp ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= input_mem_banks_bank_a_45_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1370_tmp ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= input_mem_banks_bank_a_46_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1372_tmp ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= input_mem_banks_bank_a_47_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1374_tmp ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= input_mem_banks_bank_a_48_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1376_tmp ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= input_mem_banks_bank_a_49_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1378_tmp ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= input_mem_banks_bank_a_50_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1380_tmp ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= input_mem_banks_bank_a_51_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1382_tmp ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= input_mem_banks_bank_a_52_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1384_tmp ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= input_mem_banks_bank_a_53_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1386_tmp ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= input_mem_banks_bank_a_54_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1388_tmp ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= input_mem_banks_bank_a_55_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1390_tmp ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= input_mem_banks_bank_a_56_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1392_tmp ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= input_mem_banks_bank_a_57_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1394_tmp ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= input_mem_banks_bank_a_58_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1396_tmp ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= input_mem_banks_bank_a_59_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1398_tmp ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= input_mem_banks_bank_a_60_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1400_tmp ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= input_mem_banks_bank_a_61_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1402_tmp ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= input_mem_banks_bank_a_62_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1404_tmp ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= input_mem_banks_bank_a_63_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1406_tmp ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= input_mem_banks_bank_a_64_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1408_tmp ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= input_mem_banks_bank_a_65_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1410_tmp ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= input_mem_banks_bank_a_66_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1412_tmp ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= input_mem_banks_bank_a_67_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1414_tmp ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= input_mem_banks_bank_a_68_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1416_tmp ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= input_mem_banks_bank_a_69_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1418_tmp ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= input_mem_banks_bank_a_70_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1420_tmp ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= input_mem_banks_bank_a_71_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1422_tmp ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= input_mem_banks_bank_a_72_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1424_tmp ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= input_mem_banks_bank_a_73_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1426_tmp ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= input_mem_banks_bank_a_74_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1428_tmp ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= input_mem_banks_bank_a_75_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1430_tmp ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= input_mem_banks_bank_a_76_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1432_tmp ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= input_mem_banks_bank_a_77_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1434_tmp ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= input_mem_banks_bank_a_78_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1436_tmp ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= input_mem_banks_bank_a_79_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1438_tmp ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= input_mem_banks_bank_a_80_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1440_tmp ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= input_mem_banks_bank_a_81_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1442_tmp ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= input_mem_banks_bank_a_82_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1444_tmp ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= input_mem_banks_bank_a_83_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1446_tmp ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= input_mem_banks_bank_a_84_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1448_tmp ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= input_mem_banks_bank_a_85_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1450_tmp ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= input_mem_banks_bank_a_86_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1452_tmp ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= input_mem_banks_bank_a_87_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1454_tmp ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= input_mem_banks_bank_a_88_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1456_tmp ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= input_mem_banks_bank_a_89_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1458_tmp ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= input_mem_banks_bank_a_90_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1460_tmp ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= input_mem_banks_bank_a_91_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1462_tmp ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= input_mem_banks_bank_a_92_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1464_tmp ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= input_mem_banks_bank_a_93_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1466_tmp ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= input_mem_banks_bank_a_94_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1468_tmp ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= input_mem_banks_bank_a_95_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1470_tmp ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= input_mem_banks_bank_a_96_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1472_tmp ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= input_mem_banks_bank_a_97_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1474_tmp ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= input_mem_banks_bank_a_98_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1476_tmp ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= input_mem_banks_bank_a_99_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1478_tmp ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= input_mem_banks_bank_a_100_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1480_tmp ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= input_mem_banks_bank_a_101_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1482_tmp ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= input_mem_banks_bank_a_102_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1484_tmp ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= input_mem_banks_bank_a_103_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1486_tmp ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= input_mem_banks_bank_a_104_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1488_tmp ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= input_mem_banks_bank_a_105_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1490_tmp ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= input_mem_banks_bank_a_106_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1492_tmp ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= input_mem_banks_bank_a_107_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1494_tmp ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= input_mem_banks_bank_a_108_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1496_tmp ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= input_mem_banks_bank_a_109_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1498_tmp ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= input_mem_banks_bank_a_110_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1500_tmp ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= input_mem_banks_bank_a_111_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1502_tmp ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= input_mem_banks_bank_a_112_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1504_tmp ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= input_mem_banks_bank_a_113_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1506_tmp ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= input_mem_banks_bank_a_114_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1508_tmp ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= input_mem_banks_bank_a_115_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1510_tmp ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= input_mem_banks_bank_a_116_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1512_tmp ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= input_mem_banks_bank_a_117_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1514_tmp ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= input_mem_banks_bank_a_118_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1516_tmp ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= input_mem_banks_bank_a_119_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1518_tmp ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= input_mem_banks_bank_a_120_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1520_tmp ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= input_mem_banks_bank_a_121_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1522_tmp ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= input_mem_banks_bank_a_122_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1524_tmp ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= input_mem_banks_bank_a_123_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1526_tmp ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= input_mem_banks_bank_a_124_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1528_tmp ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= input_mem_banks_bank_a_125_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1530_tmp ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= input_mem_banks_bank_a_126_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1532_tmp ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= input_mem_banks_bank_a_127_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1534_tmp ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= input_mem_banks_bank_a_128_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1536_tmp ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= input_mem_banks_bank_a_129_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1538_tmp ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= input_mem_banks_bank_a_130_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1540_tmp ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= input_mem_banks_bank_a_131_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1542_tmp ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= input_mem_banks_bank_a_132_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1544_tmp ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= input_mem_banks_bank_a_133_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1546_tmp ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= input_mem_banks_bank_a_134_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1548_tmp ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= input_mem_banks_bank_a_135_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1550_tmp ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= input_mem_banks_bank_a_136_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1552_tmp ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= input_mem_banks_bank_a_137_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1554_tmp ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= input_mem_banks_bank_a_138_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1556_tmp ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= input_mem_banks_bank_a_139_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1558_tmp ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= input_mem_banks_bank_a_140_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1560_tmp ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= input_mem_banks_bank_a_141_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1562_tmp ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= input_mem_banks_bank_a_142_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1564_tmp ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= input_mem_banks_bank_a_143_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1566_tmp ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= input_mem_banks_bank_a_144_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1568_tmp ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= input_mem_banks_bank_a_145_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1570_tmp ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= input_mem_banks_bank_a_146_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1572_tmp ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= input_mem_banks_bank_a_147_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1574_tmp ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= input_mem_banks_bank_a_148_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1576_tmp ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= input_mem_banks_bank_a_149_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1578_tmp ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= input_mem_banks_bank_a_150_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1580_tmp ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= input_mem_banks_bank_a_151_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1582_tmp ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= input_mem_banks_bank_a_152_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1584_tmp ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= input_mem_banks_bank_a_153_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1586_tmp ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= input_mem_banks_bank_a_154_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1588_tmp ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= input_mem_banks_bank_a_155_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1590_tmp ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= input_mem_banks_bank_a_156_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1592_tmp ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= input_mem_banks_bank_a_157_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1594_tmp ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= input_mem_banks_bank_a_158_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1596_tmp ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= input_mem_banks_bank_a_159_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1598_tmp ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= input_mem_banks_bank_a_160_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1600_tmp ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= input_mem_banks_bank_a_161_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1602_tmp ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= input_mem_banks_bank_a_162_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1604_tmp ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= input_mem_banks_bank_a_163_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1606_tmp ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= input_mem_banks_bank_a_164_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1608_tmp ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= input_mem_banks_bank_a_165_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1610_tmp ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= input_mem_banks_bank_a_166_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1612_tmp ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= input_mem_banks_bank_a_167_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1614_tmp ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= input_mem_banks_bank_a_168_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1616_tmp ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= input_mem_banks_bank_a_169_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1618_tmp ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= input_mem_banks_bank_a_170_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1620_tmp ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= input_mem_banks_bank_a_171_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1622_tmp ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= input_mem_banks_bank_a_172_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1624_tmp ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= input_mem_banks_bank_a_173_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1626_tmp ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= input_mem_banks_bank_a_174_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1628_tmp ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= input_mem_banks_bank_a_175_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1630_tmp ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= input_mem_banks_bank_a_176_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1632_tmp ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= input_mem_banks_bank_a_177_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1634_tmp ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= input_mem_banks_bank_a_178_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1636_tmp ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= input_mem_banks_bank_a_179_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1638_tmp ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= input_mem_banks_bank_a_180_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1640_tmp ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= input_mem_banks_bank_a_181_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1642_tmp ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= input_mem_banks_bank_a_182_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1644_tmp ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= input_mem_banks_bank_a_183_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1646_tmp ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= input_mem_banks_bank_a_184_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1648_tmp ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= input_mem_banks_bank_a_185_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1650_tmp ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= input_mem_banks_bank_a_186_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1652_tmp ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= input_mem_banks_bank_a_187_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1654_tmp ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= input_mem_banks_bank_a_188_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1656_tmp ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= input_mem_banks_bank_a_189_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1658_tmp ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= input_mem_banks_bank_a_190_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1660_tmp ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= input_mem_banks_bank_a_191_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1662_tmp ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= input_mem_banks_bank_a_192_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1664_tmp ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= input_mem_banks_bank_a_193_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1666_tmp ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= input_mem_banks_bank_a_194_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1668_tmp ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= input_mem_banks_bank_a_195_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1670_tmp ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= input_mem_banks_bank_a_196_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1672_tmp ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= input_mem_banks_bank_a_197_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1674_tmp ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= input_mem_banks_bank_a_198_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1676_tmp ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= input_mem_banks_bank_a_199_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1678_tmp ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= input_mem_banks_bank_a_200_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1680_tmp ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= input_mem_banks_bank_a_201_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1682_tmp ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= input_mem_banks_bank_a_202_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1684_tmp ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= input_mem_banks_bank_a_203_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1686_tmp ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= input_mem_banks_bank_a_204_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1688_tmp ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= input_mem_banks_bank_a_205_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1690_tmp ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= input_mem_banks_bank_a_206_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1692_tmp ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= input_mem_banks_bank_a_207_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1694_tmp ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= input_mem_banks_bank_a_208_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1696_tmp ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= input_mem_banks_bank_a_209_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1698_tmp ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= input_mem_banks_bank_a_210_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1700_tmp ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= input_mem_banks_bank_a_211_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1702_tmp ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= input_mem_banks_bank_a_212_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1704_tmp ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= input_mem_banks_bank_a_213_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1706_tmp ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= input_mem_banks_bank_a_214_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1708_tmp ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= input_mem_banks_bank_a_215_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1710_tmp ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= input_mem_banks_bank_a_216_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1712_tmp ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= input_mem_banks_bank_a_217_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1714_tmp ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= input_mem_banks_bank_a_218_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1716_tmp ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= input_mem_banks_bank_a_219_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1718_tmp ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= input_mem_banks_bank_a_220_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1720_tmp ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= input_mem_banks_bank_a_221_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1722_tmp ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= input_mem_banks_bank_a_222_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1724_tmp ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= input_mem_banks_bank_a_223_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1726_tmp ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= input_mem_banks_bank_a_224_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1728_tmp ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= input_mem_banks_bank_a_225_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1730_tmp ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= input_mem_banks_bank_a_226_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1732_tmp ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= input_mem_banks_bank_a_227_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1734_tmp ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= input_mem_banks_bank_a_228_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1736_tmp ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= input_mem_banks_bank_a_229_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1738_tmp ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= input_mem_banks_bank_a_230_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1740_tmp ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= input_mem_banks_bank_a_231_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1742_tmp ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= input_mem_banks_bank_a_232_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1744_tmp ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= input_mem_banks_bank_a_233_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1746_tmp ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= input_mem_banks_bank_a_234_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1748_tmp ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= input_mem_banks_bank_a_235_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1750_tmp ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= input_mem_banks_bank_a_236_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1752_tmp ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= input_mem_banks_bank_a_237_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1754_tmp ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= input_mem_banks_bank_a_238_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1756_tmp ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= input_mem_banks_bank_a_239_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1758_tmp ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= input_mem_banks_bank_a_240_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1760_tmp ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= input_mem_banks_bank_a_241_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1762_tmp ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= input_mem_banks_bank_a_242_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1764_tmp ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= input_mem_banks_bank_a_243_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1766_tmp ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= input_mem_banks_bank_a_244_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1768_tmp ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= input_mem_banks_bank_a_245_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1770_tmp ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= input_mem_banks_bank_a_246_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1772_tmp ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= input_mem_banks_bank_a_247_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1774_tmp ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= input_mem_banks_bank_a_248_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1776_tmp ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= input_mem_banks_bank_a_249_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1778_tmp ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= input_mem_banks_bank_a_250_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1780_tmp ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= input_mem_banks_bank_a_251_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1782_tmp ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= input_mem_banks_bank_a_252_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1784_tmp ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= input_mem_banks_bank_a_253_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1786_tmp ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= input_mem_banks_bank_a_254_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1788_tmp ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= input_mem_banks_bank_a_255_sva_dfm_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= pe_manager_base_weight_slc_pe_manager_base_weight_0_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_28_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0 <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( input_read_req_valid_and_4_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_19_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_4 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_50_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_4 <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= 4'b0000;
      rva_out_reg_data_62_56_sva_dfm_4_1 <= 7'b0000000;
      rva_out_reg_data_46_40_sva_dfm_4_1_3_0 <= 4'b0000;
      rva_out_reg_data_55_48_sva_dfm_4_1_7_4 <= 4'b0000;
      rva_out_reg_data_55_48_sva_dfm_4_1_3_0 <= 4'b0000;
    end
    else if ( and_1792_cse ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= MUX1HOT_v_4_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0,
          rva_out_reg_data_35_32_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[35:32]),
          (weight_port_read_out_data_0_4_sva_dfm_3_5_0[3:0]), {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_62_56_sva_dfm_4_1 <= MUX1HOT_v_7_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0,
          rva_out_reg_data_62_56_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[62:56]),
          weight_port_read_out_data_0_7_sva_dfm_3_6_0, {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_46_40_sva_dfm_4_1_3_0 <= MUX1HOT_v_4_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0[3:0]),
          rva_out_reg_data_46_40_sva_dfm_6_mx1_3_0, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[43:40]),
          weight_port_read_out_data_0_5_sva_dfm_3_3_0, {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_55_48_sva_dfm_4_1_7_4 <= MUX1HOT_v_4_4_2((rva_out_reg_data_55_48_sva_dfm_1_5[7:4]),
          rva_out_reg_data_55_48_sva_dfm_6_mx1_7_4, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:52]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_7_4,
          {PECore_PushAxiRsp_if_asn_61 , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65
          , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_55_48_sva_dfm_4_1_3_0 <= MUX1HOT_v_4_4_2((rva_out_reg_data_55_48_sva_dfm_1_5[3:0]),
          rva_out_reg_data_55_48_sva_dfm_6_mx1_3_0, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[51:48]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_3_0,
          {PECore_PushAxiRsp_if_asn_61 , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65
          , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_3_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_35_32_sva_dfm_6 <= 4'b0000;
      rva_out_reg_data_55_48_sva_dfm_6_rsp_0 <= 4'b0000;
      rva_out_reg_data_55_48_sva_dfm_6_rsp_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_6_rsp_1 <= 4'b0000;
    end
    else if ( and_1801_cse ) begin
      rva_out_reg_data_62_56_sva_dfm_6 <= rva_out_reg_data_62_56_sva_dfm_6_mx1;
      rva_out_reg_data_35_32_sva_dfm_6 <= rva_out_reg_data_35_32_sva_dfm_6_mx1;
      rva_out_reg_data_55_48_sva_dfm_6_rsp_0 <= rva_out_reg_data_55_48_sva_dfm_6_mx1_7_4;
      rva_out_reg_data_55_48_sva_dfm_6_rsp_1 <= rva_out_reg_data_55_48_sva_dfm_6_mx1_3_0;
      rva_out_reg_data_46_40_sva_dfm_6_rsp_1 <= rva_out_reg_data_46_40_sva_dfm_6_mx1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_13_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & ((rva_in_reg_rw_sva_5 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
        & while_stage_0_7) | PECore_PushAxiRsp_mux_13_itm_1_mx0c1) ) begin
      PECore_PushAxiRsp_mux_13_itm_1 <= MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
          weight_port_read_out_data_mux_71_nl, PECore_PushAxiRsp_mux_13_itm_1_mx0c1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ rva_in_reg_rw_sva_5) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
        & while_stage_0_7 & fsm_output ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          (weight_port_read_out_data_0_5_sva_dfm_3_7_4[3]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_5 <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_61_cse ) begin
      rva_out_reg_data_55_48_sva_dfm_1_5 <= MUX_v_8_2_2(rva_out_reg_data_55_48_sva_dfm_1_4,
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7
          <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm[7];
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0
          <= MUX_v_7_2_2(rva_out_reg_data_62_56_sva_dfm_1_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm[6:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_29_tmp ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= MUX1HOT_v_64_3_2(input_mem_banks_read_1_read_data_lpi_1_dfm_1_3,
          weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d, weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1,
          {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          , and_639_nl , nor_418_nl});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_base_input_and_tmp ) begin
      pe_manager_base_input_sva <= MUX_v_15_2_2(pe_manager_base_input_sva_dfm_3_1,
          while_if_while_if_and_2_nl, and_dcpl_240);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( (~((~((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6:4]!=3'b000)))
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9:7]!=3'b000))) & nor_718_cse
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:12]!=3'b000))) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]))
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & rva_in_PopNB_mioi_return_rsc_z_mxwt
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]==2'b00) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt))
        & while_stage_0_3)) & rva_in_reg_rw_and_6_cse ) begin
      pe_manager_base_input_sva_dfm_3_1 <= MUX_v_15_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[62:48]),
          pe_manager_base_input_sva_mx2, or_492_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_90_nl) & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_20_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_23_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_23_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_93_nl) & while_stage_0_5 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= MUX_s_1_2_2((pe_manager_base_weight_sva[0]), PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_95_nl & while_stage_0_5 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= MUX_s_1_2_2((pe_manager_base_weight_sva[0]), PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_27_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_107_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= rva_out_reg_data_30_25_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_108_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= rva_out_reg_data_23_17_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_109_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= rva_out_reg_data_15_9_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_110_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= rva_out_reg_data_35_32_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_111_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= rva_out_reg_data_39_36_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_112_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= rva_out_reg_data_46_40_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_113_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_4 <= rva_out_reg_data_62_56_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_114_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_4 <= rva_out_reg_data_55_48_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_28_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(reg_rva_in_reg_rw_sva_2_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= MUX_s_1_2_2((pe_manager_base_weight_sva_mx1_3_0[1]), PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ reg_rva_in_reg_rw_sva_2_cse) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= input_read_req_valid_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_31_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= 6'b000000;
      rva_out_reg_data_23_17_sva_dfm_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_70_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= MUX_v_6_2_2(6'b000000, (pe_manager_base_weight_sva_mx2[14:9]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
      rva_out_reg_data_23_17_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_base_weight_sva_mx2[7:1]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_115_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= rva_out_reg_data_15_9_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_116_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= rva_out_reg_data_35_32_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_117_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= rva_out_reg_data_39_36_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_118_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= rva_out_reg_data_46_40_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_119_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_3 <= rva_out_reg_data_62_56_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_120_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_3 <= rva_out_reg_data_55_48_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_33_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= 1'b0;
      input_read_req_valid_lpi_1_dfm_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
      input_read_req_valid_lpi_1_dfm_1_2 <= input_read_req_valid_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_35_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_78_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= rva_out_reg_data_15_9_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_121_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= rva_out_reg_data_35_32_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_122_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= rva_out_reg_data_39_36_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_123_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= rva_out_reg_data_46_40_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_124_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_2 <= rva_out_reg_data_62_56_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_125_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_2 <= rva_out_reg_data_55_48_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (and_dcpl_434 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        & while_stage_0_3 ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_2_1,
          PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_434 & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1==4'b0100)
        & and_dcpl_441 & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3))
        & and_dcpl_194 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_38_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_1 <= 7'b0000000;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_6_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1);
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_3;
      rva_out_reg_data_15_9_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_num_input_sva[7:1]),
          and_301_cse);
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_43_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= pe_config_is_cluster_sva;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1 <= pe_config_is_bias_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_sva_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_30_tmp ) begin
      input_mem_banks_read_read_data_sva_1 <= MUX_v_64_256_2(input_mem_banks_bank_a_mux_1_nl,
          input_mem_banks_bank_a_mux_3_nl, input_mem_banks_bank_a_mux_5_nl, input_mem_banks_bank_a_mux_7_nl,
          input_mem_banks_bank_a_mux_9_nl, input_mem_banks_bank_a_mux_11_nl, input_mem_banks_bank_a_mux_13_nl,
          input_mem_banks_bank_a_mux_15_nl, input_mem_banks_bank_a_mux_17_nl, input_mem_banks_bank_a_mux_19_nl,
          input_mem_banks_bank_a_mux_21_nl, input_mem_banks_bank_a_mux_23_nl, input_mem_banks_bank_a_mux_25_nl,
          input_mem_banks_bank_a_mux_27_nl, input_mem_banks_bank_a_mux_29_nl, input_mem_banks_bank_a_mux_31_nl,
          input_mem_banks_bank_a_mux_33_nl, input_mem_banks_bank_a_mux_35_nl, input_mem_banks_bank_a_mux_37_nl,
          input_mem_banks_bank_a_mux_39_nl, input_mem_banks_bank_a_mux_41_nl, input_mem_banks_bank_a_mux_43_nl,
          input_mem_banks_bank_a_mux_45_nl, input_mem_banks_bank_a_mux_47_nl, input_mem_banks_bank_a_mux_49_nl,
          input_mem_banks_bank_a_mux_51_nl, input_mem_banks_bank_a_mux_53_nl, input_mem_banks_bank_a_mux_55_nl,
          input_mem_banks_bank_a_mux_57_nl, input_mem_banks_bank_a_mux_59_nl, input_mem_banks_bank_a_mux_61_nl,
          input_mem_banks_bank_a_mux_63_nl, input_mem_banks_bank_a_mux_65_nl, input_mem_banks_bank_a_mux_67_nl,
          input_mem_banks_bank_a_mux_69_nl, input_mem_banks_bank_a_mux_71_nl, input_mem_banks_bank_a_mux_73_nl,
          input_mem_banks_bank_a_mux_75_nl, input_mem_banks_bank_a_mux_77_nl, input_mem_banks_bank_a_mux_79_nl,
          input_mem_banks_bank_a_mux_81_nl, input_mem_banks_bank_a_mux_83_nl, input_mem_banks_bank_a_mux_85_nl,
          input_mem_banks_bank_a_mux_87_nl, input_mem_banks_bank_a_mux_89_nl, input_mem_banks_bank_a_mux_91_nl,
          input_mem_banks_bank_a_mux_93_nl, input_mem_banks_bank_a_mux_95_nl, input_mem_banks_bank_a_mux_97_nl,
          input_mem_banks_bank_a_mux_99_nl, input_mem_banks_bank_a_mux_101_nl, input_mem_banks_bank_a_mux_103_nl,
          input_mem_banks_bank_a_mux_105_nl, input_mem_banks_bank_a_mux_107_nl, input_mem_banks_bank_a_mux_109_nl,
          input_mem_banks_bank_a_mux_111_nl, input_mem_banks_bank_a_mux_113_nl, input_mem_banks_bank_a_mux_115_nl,
          input_mem_banks_bank_a_mux_117_nl, input_mem_banks_bank_a_mux_119_nl, input_mem_banks_bank_a_mux_121_nl,
          input_mem_banks_bank_a_mux_123_nl, input_mem_banks_bank_a_mux_125_nl, input_mem_banks_bank_a_mux_127_nl,
          input_mem_banks_bank_a_mux_129_nl, input_mem_banks_bank_a_mux_131_nl, input_mem_banks_bank_a_mux_133_nl,
          input_mem_banks_bank_a_mux_135_nl, input_mem_banks_bank_a_mux_137_nl, input_mem_banks_bank_a_mux_139_nl,
          input_mem_banks_bank_a_mux_141_nl, input_mem_banks_bank_a_mux_143_nl, input_mem_banks_bank_a_mux_145_nl,
          input_mem_banks_bank_a_mux_147_nl, input_mem_banks_bank_a_mux_149_nl, input_mem_banks_bank_a_mux_151_nl,
          input_mem_banks_bank_a_mux_153_nl, input_mem_banks_bank_a_mux_155_nl, input_mem_banks_bank_a_mux_157_nl,
          input_mem_banks_bank_a_mux_159_nl, input_mem_banks_bank_a_mux_161_nl, input_mem_banks_bank_a_mux_163_nl,
          input_mem_banks_bank_a_mux_165_nl, input_mem_banks_bank_a_mux_167_nl, input_mem_banks_bank_a_mux_169_nl,
          input_mem_banks_bank_a_mux_171_nl, input_mem_banks_bank_a_mux_173_nl, input_mem_banks_bank_a_mux_175_nl,
          input_mem_banks_bank_a_mux_177_nl, input_mem_banks_bank_a_mux_179_nl, input_mem_banks_bank_a_mux_181_nl,
          input_mem_banks_bank_a_mux_183_nl, input_mem_banks_bank_a_mux_185_nl, input_mem_banks_bank_a_mux_187_nl,
          input_mem_banks_bank_a_mux_189_nl, input_mem_banks_bank_a_mux_191_nl, input_mem_banks_bank_a_mux_193_nl,
          input_mem_banks_bank_a_mux_195_nl, input_mem_banks_bank_a_mux_197_nl, input_mem_banks_bank_a_mux_199_nl,
          input_mem_banks_bank_a_mux_201_nl, input_mem_banks_bank_a_mux_203_nl, input_mem_banks_bank_a_mux_205_nl,
          input_mem_banks_bank_a_mux_207_nl, input_mem_banks_bank_a_mux_209_nl, input_mem_banks_bank_a_mux_211_nl,
          input_mem_banks_bank_a_mux_213_nl, input_mem_banks_bank_a_mux_215_nl, input_mem_banks_bank_a_mux_217_nl,
          input_mem_banks_bank_a_mux_219_nl, input_mem_banks_bank_a_mux_221_nl, input_mem_banks_bank_a_mux_223_nl,
          input_mem_banks_bank_a_mux_225_nl, input_mem_banks_bank_a_mux_227_nl, input_mem_banks_bank_a_mux_229_nl,
          input_mem_banks_bank_a_mux_231_nl, input_mem_banks_bank_a_mux_233_nl, input_mem_banks_bank_a_mux_235_nl,
          input_mem_banks_bank_a_mux_237_nl, input_mem_banks_bank_a_mux_239_nl, input_mem_banks_bank_a_mux_241_nl,
          input_mem_banks_bank_a_mux_243_nl, input_mem_banks_bank_a_mux_245_nl, input_mem_banks_bank_a_mux_247_nl,
          input_mem_banks_bank_a_mux_249_nl, input_mem_banks_bank_a_mux_251_nl, input_mem_banks_bank_a_mux_253_nl,
          input_mem_banks_bank_a_mux_255_nl, input_mem_banks_bank_a_mux_257_nl, input_mem_banks_bank_a_mux_259_nl,
          input_mem_banks_bank_a_mux_261_nl, input_mem_banks_bank_a_mux_263_nl, input_mem_banks_bank_a_mux_265_nl,
          input_mem_banks_bank_a_mux_267_nl, input_mem_banks_bank_a_mux_269_nl, input_mem_banks_bank_a_mux_271_nl,
          input_mem_banks_bank_a_mux_273_nl, input_mem_banks_bank_a_mux_275_nl, input_mem_banks_bank_a_mux_277_nl,
          input_mem_banks_bank_a_mux_279_nl, input_mem_banks_bank_a_mux_281_nl, input_mem_banks_bank_a_mux_283_nl,
          input_mem_banks_bank_a_mux_285_nl, input_mem_banks_bank_a_mux_287_nl, input_mem_banks_bank_a_mux_289_nl,
          input_mem_banks_bank_a_mux_291_nl, input_mem_banks_bank_a_mux_293_nl, input_mem_banks_bank_a_mux_295_nl,
          input_mem_banks_bank_a_mux_297_nl, input_mem_banks_bank_a_mux_299_nl, input_mem_banks_bank_a_mux_301_nl,
          input_mem_banks_bank_a_mux_303_nl, input_mem_banks_bank_a_mux_305_nl, input_mem_banks_bank_a_mux_307_nl,
          input_mem_banks_bank_a_mux_309_nl, input_mem_banks_bank_a_mux_311_nl, input_mem_banks_bank_a_mux_313_nl,
          input_mem_banks_bank_a_mux_315_nl, input_mem_banks_bank_a_mux_317_nl, input_mem_banks_bank_a_mux_319_nl,
          input_mem_banks_bank_a_mux_321_nl, input_mem_banks_bank_a_mux_323_nl, input_mem_banks_bank_a_mux_325_nl,
          input_mem_banks_bank_a_mux_327_nl, input_mem_banks_bank_a_mux_329_nl, input_mem_banks_bank_a_mux_331_nl,
          input_mem_banks_bank_a_mux_333_nl, input_mem_banks_bank_a_mux_335_nl, input_mem_banks_bank_a_mux_337_nl,
          input_mem_banks_bank_a_mux_339_nl, input_mem_banks_bank_a_mux_341_nl, input_mem_banks_bank_a_mux_343_nl,
          input_mem_banks_bank_a_mux_345_nl, input_mem_banks_bank_a_mux_347_nl, input_mem_banks_bank_a_mux_349_nl,
          input_mem_banks_bank_a_mux_351_nl, input_mem_banks_bank_a_mux_353_nl, input_mem_banks_bank_a_mux_355_nl,
          input_mem_banks_bank_a_mux_357_nl, input_mem_banks_bank_a_mux_359_nl, input_mem_banks_bank_a_mux_361_nl,
          input_mem_banks_bank_a_mux_363_nl, input_mem_banks_bank_a_mux_365_nl, input_mem_banks_bank_a_mux_367_nl,
          input_mem_banks_bank_a_mux_369_nl, input_mem_banks_bank_a_mux_371_nl, input_mem_banks_bank_a_mux_373_nl,
          input_mem_banks_bank_a_mux_375_nl, input_mem_banks_bank_a_mux_377_nl, input_mem_banks_bank_a_mux_379_nl,
          input_mem_banks_bank_a_mux_381_nl, input_mem_banks_bank_a_mux_383_nl, input_mem_banks_bank_a_mux_385_nl,
          input_mem_banks_bank_a_mux_387_nl, input_mem_banks_bank_a_mux_389_nl, input_mem_banks_bank_a_mux_391_nl,
          input_mem_banks_bank_a_mux_393_nl, input_mem_banks_bank_a_mux_395_nl, input_mem_banks_bank_a_mux_397_nl,
          input_mem_banks_bank_a_mux_399_nl, input_mem_banks_bank_a_mux_401_nl, input_mem_banks_bank_a_mux_403_nl,
          input_mem_banks_bank_a_mux_405_nl, input_mem_banks_bank_a_mux_407_nl, input_mem_banks_bank_a_mux_409_nl,
          input_mem_banks_bank_a_mux_411_nl, input_mem_banks_bank_a_mux_413_nl, input_mem_banks_bank_a_mux_415_nl,
          input_mem_banks_bank_a_mux_417_nl, input_mem_banks_bank_a_mux_419_nl, input_mem_banks_bank_a_mux_421_nl,
          input_mem_banks_bank_a_mux_423_nl, input_mem_banks_bank_a_mux_425_nl, input_mem_banks_bank_a_mux_427_nl,
          input_mem_banks_bank_a_mux_429_nl, input_mem_banks_bank_a_mux_431_nl, input_mem_banks_bank_a_mux_433_nl,
          input_mem_banks_bank_a_mux_435_nl, input_mem_banks_bank_a_mux_437_nl, input_mem_banks_bank_a_mux_439_nl,
          input_mem_banks_bank_a_mux_441_nl, input_mem_banks_bank_a_mux_443_nl, input_mem_banks_bank_a_mux_445_nl,
          input_mem_banks_bank_a_mux_447_nl, input_mem_banks_bank_a_mux_449_nl, input_mem_banks_bank_a_mux_451_nl,
          input_mem_banks_bank_a_mux_453_nl, input_mem_banks_bank_a_mux_455_nl, input_mem_banks_bank_a_mux_457_nl,
          input_mem_banks_bank_a_mux_459_nl, input_mem_banks_bank_a_mux_461_nl, input_mem_banks_bank_a_mux_463_nl,
          input_mem_banks_bank_a_mux_465_nl, input_mem_banks_bank_a_mux_467_nl, input_mem_banks_bank_a_mux_469_nl,
          input_mem_banks_bank_a_mux_471_nl, input_mem_banks_bank_a_mux_473_nl, input_mem_banks_bank_a_mux_475_nl,
          input_mem_banks_bank_a_mux_477_nl, input_mem_banks_bank_a_mux_479_nl, input_mem_banks_bank_a_mux_481_nl,
          input_mem_banks_bank_a_mux_483_nl, input_mem_banks_bank_a_mux_485_nl, input_mem_banks_bank_a_mux_487_nl,
          input_mem_banks_bank_a_mux_489_nl, input_mem_banks_bank_a_mux_491_nl, input_mem_banks_bank_a_mux_493_nl,
          input_mem_banks_bank_a_mux_495_nl, input_mem_banks_bank_a_mux_497_nl, input_mem_banks_bank_a_mux_499_nl,
          input_mem_banks_bank_a_mux_501_nl, input_mem_banks_bank_a_mux_503_nl, input_mem_banks_bank_a_mux_505_nl,
          input_mem_banks_bank_a_mux_507_nl, input_mem_banks_bank_a_mux_509_nl, input_mem_banks_bank_a_mux_511_nl,
          rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_39_36_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_1_1 <= 7'b0000000;
      rva_out_reg_data_62_56_sva_dfm_1_1 <= 7'b0000000;
      rva_out_reg_data_55_48_sva_dfm_1_1 <= 8'b00000000;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_85_cse ) begin
      rva_out_reg_data_35_32_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl
          & (signext_4_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1)) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_39_36_sva_dfm_1_1 <= (pe_manager_base_bias_sva[7:4]) & ({{3{and_301_cse}},
          and_301_cse}) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_46_40_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl
          & (signext_7_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1)) & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_62_56_sva_dfm_1_1 <= (pe_manager_base_input_sva_mx2[14:8])
          & ({{6{and_301_cse}}, and_301_cse}) & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_55_48_sva_dfm_1_1 <= pe_manager_base_input_sva_mx1_7_0 & ({{7{and_301_cse}},
          and_301_cse}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1_1 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_5_mux_17_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_17_itm_1_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_17_itm_1_5_0 <= 6'b000000;
    end
    else if ( weight_mem_run_3_for_5_and_222_ssc ) begin
      weight_mem_run_3_for_5_mux_17_itm_1_7 <= MUX1HOT_s_1_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006[7]),
          (weight_port_read_out_data_2_1_sva_dfm_1[7]), weight_port_read_out_data_0_2_sva_dfm_mx0w2_7,
          {and_536_itm , nor_413_itm , while_and_24_cse});
      weight_mem_run_3_for_5_mux_17_itm_1_6 <= MUX1HOT_s_1_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006[6]),
          (weight_port_read_out_data_2_1_sva_dfm_1[6]), weight_port_read_out_data_0_2_sva_dfm_mx0w2_6,
          (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0[6]),
          {and_536_itm , nor_413_itm , while_and_24_cse , while_and_23_cse});
      weight_mem_run_3_for_5_mux_17_itm_1_5_0 <= MUX1HOT_v_6_4_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006[5:0]),
          (weight_port_read_out_data_2_1_sva_dfm_1[5:0]), weight_port_read_out_data_0_2_sva_dfm_mx0w2_5_0,
          (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0[5:0]),
          {and_536_itm , nor_413_itm , while_and_24_cse , while_and_23_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7_4
          <= 4'b0000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0
          <= 4'b0000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_1_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7_4
          <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm[7:4];
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0
          <= MUX_v_4_2_2(rva_out_reg_data_39_36_sva_dfm_1_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm[3:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0
          <= 7'b0000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4
          <= 4'b0000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0
          <= 4'b0000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_7_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_8_nl & (~ or_dcpl_297);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_38_nl,
          not_2208_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4
          <= MUX_v_4_2_2(4'b0000, weight_mem_banks_load_store_for_else_mux1h_15_nl,
          not_2209_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0
          <= MUX_v_4_2_2(4'b0000, weight_mem_banks_load_store_for_else_mux1h_39_nl,
          not_2210_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6
          <= 2'b00;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0
          <= 6'b000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0
          <= 7'b0000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_17_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6
          <= MUX_v_2_2_2(2'b00, weight_mem_banks_load_store_for_else_mux1h_22_nl,
          not_2211_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0
          <= MUX_v_6_2_2(6'b000000, weight_mem_banks_load_store_for_else_mux1h_40_nl,
          not_2212_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_27_nl & (~ or_dcpl_297);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_41_nl,
          not_2214_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_32_nl & (~ or_dcpl_297);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_42_nl,
          not_2216_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_1_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_1_rsp_0 <= 3'b000;
    end
    else if ( weight_port_read_out_data_and_86_cse ) begin
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_2_sva_dfm_2_7;
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_3_sva_dfm_2_7;
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_0_sva_dfm_2_7_1;
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_1_sva_dfm_2_7_1;
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_1_rsp_0 <= weight_port_read_out_data_0_2_sva_dfm_2_6_1;
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_1_rsp_0 <= weight_port_read_out_data_0_3_sva_dfm_2_6_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_2_7_1 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_2_7_1 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_2_6_1 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_2_6_4_1 <= 3'b000;
    end
    else if ( weight_port_read_out_data_and_90_ssc ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_7 <= weight_mem_run_3_for_5_mux_17_itm_1_7;
      weight_port_read_out_data_0_3_sva_dfm_2_7 <= weight_port_read_out_data_0_3_sva_dfm_1_7;
      weight_port_read_out_data_0_0_sva_dfm_2_7_1 <= input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_7;
      weight_port_read_out_data_0_1_sva_dfm_2_7_1 <= input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_7;
      weight_port_read_out_data_0_2_sva_dfm_2_6_1 <= weight_mem_run_3_for_5_mux_17_itm_1_6;
      weight_port_read_out_data_0_3_sva_dfm_2_6_4_1 <= weight_port_read_out_data_0_3_sva_dfm_1_6_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_7 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_1_6_4 <= 3'b000;
      weight_port_read_out_data_0_3_sva_dfm_1_3_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_94_ssc ) begin
      weight_port_read_out_data_0_3_sva_dfm_1_7 <= weight_port_read_out_data_0_3_sva_dfm_mx0w0_7;
      weight_port_read_out_data_0_3_sva_dfm_1_6_4 <= MUX_v_3_2_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0[6:4]),
          weight_port_read_out_data_0_3_sva_dfm_mx0w0_6_4, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
      weight_port_read_out_data_0_3_sva_dfm_1_3_0 <= MUX_v_4_2_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0[3:0]),
          weight_port_read_out_data_0_3_sva_dfm_mx0w0_3_0, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_7
          <= 1'b0;
      input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_6_0
          <= 7'b0000000;
      input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_7
          <= 1'b0;
      input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_ssc ) begin
      input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_7
          <= MUX_s_1_2_2((input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[7]), weight_port_read_out_data_0_1_sva_dfm_mx0w1_7,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
      input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_6_0
          <= MUX_v_7_2_2((input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[6:0]), weight_port_read_out_data_0_1_sva_dfm_mx0w1_6_0,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
      input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_7
          <= MUX_s_1_2_2((input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[15]), weight_port_read_out_data_0_0_sva_dfm_mx0w1_7,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
      input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_6_0
          <= MUX_v_7_2_2((input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[14:8]),
          weight_port_read_out_data_0_0_sva_dfm_mx0w1_6_0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_6_sva_dfm_2_7_4 <= 4'b0000;
      weight_port_read_out_data_0_6_sva_dfm_2_3_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_1_ssc ) begin
      weight_port_read_out_data_0_6_sva_dfm_2_7_4 <= MUX_v_4_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000[7:4]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_7_4,
          while_and_24_cse);
      weight_port_read_out_data_0_6_sva_dfm_2_3_0 <= MUX_v_4_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000[3:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_3_0,
          while_and_24_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_7_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_4_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_4_sva_dfm_2_6 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_2_7_1 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_2_6_4 <= 3'b000;
      weight_port_read_out_data_0_2_sva_dfm_2_7_1 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_2_6 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_2_7 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_56_cse ) begin
      weight_port_read_out_data_0_7_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_7_sva_dfm_3_7,
          Datapath_for_4_ProductSum_for_acc_5_cmp_8_a_mx1_7, and_dcpl_375);
      weight_port_read_out_data_0_4_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_4_sva_dfm_3_7,
          Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_7, and_dcpl_375);
      weight_port_read_out_data_0_4_sva_dfm_2_6 <= MUX_s_1_2_2(weight_port_read_out_data_0_4_sva_dfm_3_6,
          Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_6, and_dcpl_375);
      weight_port_read_out_data_0_3_sva_dfm_2_7_1 <= MUX_s_1_2_2(weight_port_read_out_data_0_3_sva_dfm_mx0w0_7,
          Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_7, and_dcpl_375);
      weight_port_read_out_data_0_3_sva_dfm_2_6_4 <= MUX_v_3_2_2(weight_port_read_out_data_0_3_sva_dfm_mx0w0_6_4,
          Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_6_4, and_dcpl_375);
      weight_port_read_out_data_0_2_sva_dfm_2_7_1 <= MUX_s_1_2_2(weight_port_read_out_data_0_2_sva_dfm_mx0w2_7,
          Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_7, and_dcpl_375);
      weight_port_read_out_data_0_2_sva_dfm_2_6 <= MUX_s_1_2_2(weight_port_read_out_data_0_2_sva_dfm_mx0w2_6,
          Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_6, and_dcpl_375);
      weight_port_read_out_data_0_1_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_1_sva_dfm_mx0w1_7,
          Datapath_for_4_ProductSum_for_acc_5_cmp_5_a_mx1_7, and_dcpl_375);
      weight_port_read_out_data_0_0_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w1_7,
          weight_port_read_out_data_0_0_sva_dfm_3_7, and_dcpl_375);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_7_sva_dfm_2_6_0 <= 7'b0000000;
    end
    else if ( mux_887_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_7_sva_dfm_2_6_0 <= MUX_v_7_2_2(weight_port_read_out_data_0_7_sva_dfm_3_6_0,
          Datapath_for_4_ProductSum_for_acc_5_cmp_8_a_mx1_6_0, and_dcpl_375);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_5_sva_dfm_2_7_4 <= 4'b0000;
      weight_port_read_out_data_0_5_sva_dfm_2_3_0 <= 4'b0000;
    end
    else if ( and_1835_cse ) begin
      weight_port_read_out_data_0_5_sva_dfm_2_7_4 <= MUX_v_4_2_2(weight_port_read_out_data_0_5_sva_dfm_3_7_4,
          Datapath_for_4_ProductSum_for_acc_5_cmp_7_a_mx1_7_4, and_dcpl_375);
      weight_port_read_out_data_0_5_sva_dfm_2_3_0 <= MUX_v_4_2_2(weight_port_read_out_data_0_5_sva_dfm_3_3_0,
          Datapath_for_4_ProductSum_for_acc_5_cmp_7_a_mx1_3_0, and_dcpl_375);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_4_sva_dfm_2_5_0 <= 6'b000000;
    end
    else if ( mux_896_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_4_sva_dfm_2_5_0 <= MUX_v_6_2_2(weight_port_read_out_data_0_4_sva_dfm_3_5_0,
          Datapath_for_4_ProductSum_for_acc_5_cmp_7_c_mx1_5_0, and_dcpl_375);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_3_0 <= 4'b0000;
    end
    else if ( mux_899_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_3_0 <= MUX_v_4_2_2(weight_port_read_out_data_0_3_sva_dfm_mx0w0_3_0,
          Datapath_for_4_ProductSum_for_acc_5_cmp_6_a_mx1_3_0, and_dcpl_375);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_5_0 <= 6'b000000;
    end
    else if ( mux_902_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_5_0 <= MUX_v_6_2_2(weight_port_read_out_data_0_2_sva_dfm_mx0w2_5_0,
          Datapath_for_4_ProductSum_for_acc_5_cmp_6_c_mx1_5_0, and_dcpl_375);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_6_0 <= 7'b0000000;
    end
    else if ( mux_905_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_6_0 <= MUX_v_7_2_2(weight_port_read_out_data_0_1_sva_dfm_mx0w1_6_0,
          Datapath_for_4_ProductSum_for_acc_5_cmp_5_a_mx1_6_0, and_dcpl_375);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0 <= 7'b0000000;
    end
    else if ( mux_908_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0 <= MUX_v_7_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w1_6_0,
          weight_port_read_out_data_0_0_sva_dfm_3_6_0, and_dcpl_375);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_99_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1 <= weight_port_read_out_data_0_0_sva_dfm_2_6_0_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_100_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_1 <= weight_port_read_out_data_0_1_sva_dfm_2_6_0_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_6_rsp_0 <= 3'b000;
      rva_out_reg_data_15_9_sva_dfm_8_rsp_0 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_34_cse ) begin
      rva_out_reg_data_23_17_sva_dfm_6_rsp_0 <= rva_out_reg_data_23_17_sva_dfm_5_6_4;
      rva_out_reg_data_15_9_sva_dfm_8_rsp_0 <= rva_out_reg_data_15_9_sva_dfm_7_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_6_rsp_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_126_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_6_rsp_1 <= rva_out_reg_data_23_17_sva_dfm_5_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_8_rsp_1 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_127_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_8_rsp_1 <= rva_out_reg_data_15_9_sva_dfm_7_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3_rsp_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_128_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_46_40_sva_dfm_4_2_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3_rsp_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_129_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_55_48_sva_dfm_4_2_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3_rsp_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_130_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_55_48_sva_dfm_4_2_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_5_6_4 <= 3'b000;
      rva_out_reg_data_15_9_sva_dfm_7_6 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_42_cse ) begin
      rva_out_reg_data_23_17_sva_dfm_5_6_4 <= weight_port_read_out_data_0_3_sva_dfm_1_6_4;
      rva_out_reg_data_15_9_sva_dfm_7_6 <= weight_mem_run_3_for_5_mux_17_itm_1_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_5_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_131_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_5_3_0 <= weight_port_read_out_data_0_3_sva_dfm_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_7_5_0 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_132_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_7_5_0 <= weight_mem_run_3_for_5_mux_17_itm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_101_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0_1 <= input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_6_0_1 <= 7'b0000000;
    end
    else if ( weight_port_read_out_data_and_102_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_6_0_1 <= input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_133_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2_3_0 <= rva_out_reg_data_46_40_sva_dfm_4_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2_7_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_134_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2_7_4 <= rva_out_reg_data_55_48_sva_dfm_4_1_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_135_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2_3_0 <= rva_out_reg_data_55_48_sva_dfm_4_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_1_3 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_1_2 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_1_1_0 <= 2'b00;
      rva_out_reg_data_46_40_sva_dfm_4_1_6_4 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_51_cse ) begin
      rva_out_reg_data_39_36_sva_dfm_4_1_3 <= MUX1HOT_s_1_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0[3]),
          rva_out_reg_data_39_36_sva_dfm_6_mx1_3, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[39]),
          weight_port_read_out_data_0_4_sva_dfm_3_7, {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_39_36_sva_dfm_4_1_2 <= MUX1HOT_s_1_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0[2]),
          rva_out_reg_data_39_36_sva_dfm_6_mx1_2, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[38]),
          weight_port_read_out_data_0_4_sva_dfm_3_6, {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_39_36_sva_dfm_4_1_1_0 <= MUX1HOT_v_2_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0[1:0]),
          rva_out_reg_data_39_36_sva_dfm_6_mx1_1_0, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[37:36]),
          (weight_port_read_out_data_0_4_sva_dfm_3_5_0[5:4]), {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_46_40_sva_dfm_4_1_6_4 <= MUX1HOT_v_3_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0[6:4]),
          rva_out_reg_data_46_40_sva_dfm_6_mx1_6_4, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[46:44]),
          (weight_port_read_out_data_0_5_sva_dfm_3_7_4[2:0]), {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_6_rsp_0 <= 3'b000;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_0 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_1 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_2 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_56_cse ) begin
      rva_out_reg_data_46_40_sva_dfm_6_rsp_0 <= rva_out_reg_data_46_40_sva_dfm_6_mx1_6_4;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_0 <= rva_out_reg_data_39_36_sva_dfm_6_mx1_3;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_1 <= rva_out_reg_data_39_36_sva_dfm_6_mx1_2;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_2 <= rva_out_reg_data_39_36_sva_dfm_6_mx1_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_1_rsp_1 <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_103_enex5 ) begin
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_1_rsp_1 <= weight_port_read_out_data_0_2_sva_dfm_2_5_0_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_1_rsp_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_104_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_1_rsp_1 <= weight_port_read_out_data_0_3_sva_dfm_2_3_0_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_5_0_1 <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_105_enex5 ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_5_0_1 <= weight_mem_run_3_for_5_mux_17_itm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_3_0_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_106_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_3_0_1 <= weight_port_read_out_data_0_3_sva_dfm_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_10_6 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_8_6_4 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_14_cse ) begin
      rva_out_reg_data_15_9_sva_dfm_10_6 <= reg_rva_out_reg_data_15_9_sva_dfm_9_ftd;
      rva_out_reg_data_23_17_sva_dfm_8_6_4 <= reg_rva_out_reg_data_23_17_sva_dfm_7_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_10_5_0 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_136_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_10_5_0 <= reg_rva_out_reg_data_15_9_sva_dfm_9_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_8_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_137_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_8_3_0 <= reg_rva_out_reg_data_23_17_sva_dfm_7_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_5_7_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_138_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_5_7_4 <= reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_5_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_139_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_5_3_0 <= reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_5_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_140_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_5_3_0 <= reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_5_0 <=
          6'b000000;
    end
    else if ( weight_port_read_out_data_and_107_enex5 ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_2_5_0 <=
          reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_5_0 <=
          6'b000000;
    end
    else if ( weight_port_read_out_data_and_108_enex5 ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_2_5_0 <=
          reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_5_0_rsp_1
          <= 5'b00000;
    end
    else if ( weight_port_read_out_data_and_109_enex5 ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_2_5_0_rsp_1
          <= reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_5_6_0_rsp_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_110_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_5_6_0_rsp_1 <= reg_weight_port_read_out_data_0_3_sva_dfm_4_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_93_enex5 | rva_out_reg_data_and_90_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_7_enexo <= rva_out_reg_data_and_93_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_98_enex5 | rva_out_reg_data_and_91_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_4_enexo <= rva_out_reg_data_and_98_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_96_enex5 | rva_out_reg_data_and_92_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_4_enexo <= rva_out_reg_data_and_96_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_35_enex5 | input_mem_banks_read_read_data_and_31_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2_enexo
          <= input_mem_banks_read_read_data_and_35_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_36_enex5 | input_mem_banks_read_read_data_and_32_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2_enexo
          <= input_mem_banks_read_read_data_and_36_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_37_enex5 | input_mem_banks_read_read_data_and_33_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2_enexo
          <= input_mem_banks_read_read_data_and_37_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_38_enex5 | input_mem_banks_read_read_data_and_34_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2_enexo
          <= input_mem_banks_read_read_data_and_38_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_15_0_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1197_cse | act_port_reg_data_and_30_enex5 ) begin
      reg_act_port_reg_data_15_0_sva_dfm_1_1_enexo <= and_1197_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_239_224_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1197_cse | act_port_reg_data_and_31_enex5 ) begin
      reg_act_port_reg_data_239_224_sva_dfm_1_1_enexo <= and_1197_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_47_32_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1197_cse | act_port_reg_data_and_32_enex5 ) begin
      reg_act_port_reg_data_47_32_sva_dfm_1_1_enexo <= and_1197_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_207_192_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1197_cse | act_port_reg_data_and_33_enex5 ) begin
      reg_act_port_reg_data_207_192_sva_dfm_1_1_enexo <= and_1197_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_175_160_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1197_cse | act_port_reg_data_and_34_enex5 ) begin
      reg_act_port_reg_data_175_160_sva_dfm_1_1_enexo <= and_1197_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_111_96_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1197_cse | act_port_reg_data_and_35_enex5 ) begin
      reg_act_port_reg_data_111_96_sva_dfm_1_1_enexo <= and_1197_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_reg_data_143_128_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( and_1197_cse | act_port_reg_data_and_36_enex5 ) begin
      reg_act_port_reg_data_143_128_sva_dfm_1_1_enexo <= and_1197_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp | weight_port_read_out_data_and_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_000000
          <= data_in_tmp_operator_2_for_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 | input_mem_banks_read_1_read_data_and_2_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= input_mem_banks_read_1_read_data_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( weight_read_addrs_and_9_cse | weight_read_addrs_and_7_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= weight_read_addrs_and_9_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1_enexo <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1_enexo <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_23_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_23_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= 1'b1;
    end
    else if ( weight_read_addrs_and_9_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= weight_read_addrs_and_9_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_2_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1_enexo_1 <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1_enexo_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_23_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_23_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo_1
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0_enexo_1
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_17_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= 1'b1;
    end
    else if ( weight_read_addrs_and_9_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= weight_read_addrs_and_9_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= 1'b1;
    end
    else if ( operator_15_false_1_and_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= operator_15_false_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_32_enex5 | weight_write_data_data_and_24_enex5
        ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_32_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_33_enex5 | weight_write_data_data_and_25_enex5
        ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_33_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_34_enex5 | weight_write_data_data_and_26_enex5
        ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_34_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_35_enex5 | weight_write_data_data_and_27_enex5
        ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_35_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_36_enex5 | weight_write_data_data_and_28_enex5
        ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_36_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_37_enex5 | weight_write_data_data_and_29_enex5
        ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_37_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_38_enex5 | weight_write_data_data_and_30_enex5
        ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_38_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_39_enex5 | weight_write_data_data_and_31_enex5
        ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_39_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_write_addrs_and_2_enex5 | weight_write_addrs_and_enex5 ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= weight_write_addrs_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_32_enex5 ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_33_enex5 ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_34_enex5 ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_35_enex5 ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_36_enex5 ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_37_enex5 ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_38_enex5 ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_write_data_data_and_39_enex5 ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_input_enexo <= 1'b1;
    end
    else if ( pe_manager_base_input_and_tmp | weight_write_addrs_and_2_enex5 ) begin
      reg_pe_manager_base_input_enexo <= pe_manager_base_input_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_read_addrs_and_28_enex5 ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_config_num_output_enexo <= 1'b1;
    end
    else if ( pe_config_num_manager_and_cse | pe_config_UpdateManagerCounter_if_if_and_enex5
        ) begin
      reg_pe_config_num_output_enexo <= pe_config_num_manager_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_15_cse | weight_read_addrs_and_29_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= while_if_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_data_sva_1_enexo <= 1'b1;
    end
    else if ( rva_in_reg_data_and_tmp | PEManager_15U_PEManagerWrite_and_enex5 )
        begin
      reg_rva_in_reg_data_sva_1_enexo <= rva_in_reg_data_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_99_enex5 | weight_port_read_out_data_and_95_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_99_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_39_enex5 | input_mem_banks_read_read_data_and_35_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= input_mem_banks_read_read_data_and_39_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_100_enex5 | weight_port_read_out_data_and_96_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_3_1_enexo <= weight_port_read_out_data_and_100_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_40_enex5 | input_mem_banks_read_read_data_and_36_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo
          <= input_mem_banks_read_read_data_and_40_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_103_enex5 | weight_port_read_out_data_and_97_enex5
        ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_2_enexo <= weight_port_read_out_data_and_103_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_41_enex5 | input_mem_banks_read_read_data_and_37_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= input_mem_banks_read_read_data_and_41_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_42_enex5 | input_mem_banks_read_read_data_and_38_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= input_mem_banks_read_read_data_and_42_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_enex5 | input_mem_banks_read_1_read_data_and_3_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_1_read_data_and_4_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_101_enex5 | rva_out_reg_data_and_93_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= rva_out_reg_data_and_101_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_126_enex5 | rva_out_reg_data_and_94_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_1_enexo <= rva_out_reg_data_and_126_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_127_enex5 | rva_out_reg_data_and_95_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_1_enexo <= rva_out_reg_data_and_127_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_104_enex5 | weight_port_read_out_data_and_98_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_2_enexo <= weight_port_read_out_data_and_104_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_102_enex5 | rva_out_reg_data_and_96_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= rva_out_reg_data_and_102_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_128_enex5 | rva_out_reg_data_and_97_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_128_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_103_enex5 | rva_out_reg_data_and_98_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo <= rva_out_reg_data_and_103_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_129_enex5 | rva_out_reg_data_and_99_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo <= rva_out_reg_data_and_129_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_130_enex5 | rva_out_reg_data_and_100_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_130_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= 1'b1;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_1_for_and_cse | weight_mem_write_arbxbar_xbar_for_empty_and_enex5
        ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= weight_mem_write_arbxbar_xbar_for_1_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_27_enex5 | input_mem_banks_read_read_data_and_39_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo <= input_mem_banks_read_read_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_27_enex5 | input_mem_banks_read_read_data_and_40_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_1 <= input_mem_banks_read_read_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_2 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_27_enex5 | input_mem_banks_read_read_data_and_41_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_2 <= input_mem_banks_read_read_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_3 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_27_enex5 | input_mem_banks_read_read_data_and_42_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_3 <= input_mem_banks_read_read_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_5_enex5 | input_mem_banks_read_1_read_data_and_4_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= input_mem_banks_read_1_read_data_and_5_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_104_enex5 | rva_out_reg_data_and_101_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= rva_out_reg_data_and_104_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_105_enex5 | rva_out_reg_data_and_102_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= rva_out_reg_data_and_105_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_106_enex5 | rva_out_reg_data_and_103_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo <= rva_out_reg_data_and_106_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_28_enex5 | input_mem_banks_read_read_data_and_27_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0_enexo <= input_mem_banks_read_read_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_189_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1656_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_189_sva_dfm_2_enexo <= and_1656_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_208_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1694_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_208_sva_dfm_2_enexo <= and_1694_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_21_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1320_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_21_sva_dfm_2_enexo <= and_1320_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_188_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1654_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_188_sva_dfm_2_enexo <= and_1654_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_22_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1322_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_22_sva_dfm_2_enexo <= and_1322_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_249_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1776_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_249_sva_dfm_2_enexo <= and_1776_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_221_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1720_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_221_sva_dfm_2_enexo <= and_1720_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_113_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1504_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_113_sva_dfm_2_enexo <= and_1504_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_88_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1454_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_88_sva_dfm_2_enexo <= and_1454_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_13_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1304_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_13_sva_dfm_2_enexo <= and_1304_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_27_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1332_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_27_sva_dfm_2_enexo <= and_1332_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_72_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1422_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_72_sva_dfm_2_enexo <= and_1422_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_46_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1370_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_46_sva_dfm_2_enexo <= and_1370_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_132_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1542_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_132_sva_dfm_2_enexo <= and_1542_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_155_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1588_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_155_sva_dfm_2_enexo <= and_1588_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_157_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1592_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_157_sva_dfm_2_enexo <= and_1592_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_243_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1764_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_243_sva_dfm_2_enexo <= and_1764_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_149_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1576_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_149_sva_dfm_2_enexo <= and_1576_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_49_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1376_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_49_sva_dfm_2_enexo <= and_1376_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_220_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1718_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_220_sva_dfm_2_enexo <= and_1718_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_90_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1458_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_90_sva_dfm_2_enexo <= and_1458_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_83_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1444_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_83_sva_dfm_2_enexo <= and_1444_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_81_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1440_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_81_sva_dfm_2_enexo <= and_1440_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_241_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1760_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_241_sva_dfm_2_enexo <= and_1760_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_50_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1378_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_50_sva_dfm_2_enexo <= and_1378_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_96_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1470_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_96_sva_dfm_2_enexo <= and_1470_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_123_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1524_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_123_sva_dfm_2_enexo <= and_1524_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_12_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1302_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_12_sva_dfm_2_enexo <= and_1302_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_250_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1778_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_250_sva_dfm_2_enexo <= and_1778_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_248_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1774_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_248_sva_dfm_2_enexo <= and_1774_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_246_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1770_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_246_sva_dfm_2_enexo <= and_1770_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_95_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1468_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_95_sva_dfm_2_enexo <= and_1468_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_255_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1788_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_255_sva_dfm_2_enexo <= and_1788_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_17_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1312_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_17_sva_dfm_2_enexo <= and_1312_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_235_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1748_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_235_sva_dfm_2_enexo <= and_1748_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_214_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1706_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_214_sva_dfm_2_enexo <= and_1706_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_251_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1780_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_251_sva_dfm_2_enexo <= and_1780_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_read_addrs_sva_1_1_enexo <= 1'b1;
    end
    else if ( PECoreRun_wen | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_read_addrs_sva_1_1_enexo <= PECoreRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_231_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1740_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_231_sva_dfm_2_enexo <= and_1740_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_104_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1486_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_104_sva_dfm_2_enexo <= and_1486_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_142_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1562_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_142_sva_dfm_2_enexo <= and_1562_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_109_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1496_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_109_sva_dfm_2_enexo <= and_1496_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_36_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1350_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_36_sva_dfm_2_enexo <= and_1350_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_8_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1294_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_8_sva_dfm_2_enexo <= and_1294_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_19_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1316_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_19_sva_dfm_2_enexo <= and_1316_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_181_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1640_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_181_sva_dfm_2_enexo <= and_1640_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_177_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1632_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_177_sva_dfm_2_enexo <= and_1632_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_191_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1660_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_191_sva_dfm_2_enexo <= and_1660_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_4_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1286_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_4_sva_dfm_2_enexo <= and_1286_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_204_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1686_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_204_sva_dfm_2_enexo <= and_1686_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_53_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1384_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_53_sva_dfm_2_enexo <= and_1384_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_116_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1510_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_116_sva_dfm_2_enexo <= and_1510_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_139_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1556_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_139_sva_dfm_2_enexo <= and_1556_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_110_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1498_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_110_sva_dfm_2_enexo <= and_1498_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_136_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1550_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_136_sva_dfm_2_enexo <= and_1550_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_91_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1460_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_91_sva_dfm_2_enexo <= and_1460_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_55_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1388_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_55_sva_dfm_2_enexo <= and_1388_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_68_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1414_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_68_sva_dfm_2_enexo <= and_1414_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_224_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1726_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_224_sva_dfm_2_enexo <= and_1726_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_223_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1724_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_223_sva_dfm_2_enexo <= and_1724_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_93_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1464_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_93_sva_dfm_2_enexo <= and_1464_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_75_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1428_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_75_sva_dfm_2_enexo <= and_1428_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_135_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1548_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_135_sva_dfm_2_enexo <= and_1548_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_150_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1578_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_150_sva_dfm_2_enexo <= and_1578_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_108_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1494_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_108_sva_dfm_2_enexo <= and_1494_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_169_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1616_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_169_sva_dfm_2_enexo <= and_1616_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_52_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1382_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_52_sva_dfm_2_enexo <= and_1382_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_240_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1758_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_240_sva_dfm_2_enexo <= and_1758_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_213_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1704_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_213_sva_dfm_2_enexo <= and_1704_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_121_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1520_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_121_sva_dfm_2_enexo <= and_1520_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_14_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1306_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_14_sva_dfm_2_enexo <= and_1306_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_192_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1662_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_192_sva_dfm_2_enexo <= and_1662_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_194_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1666_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_194_sva_dfm_2_enexo <= and_1666_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_172_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1622_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_172_sva_dfm_2_enexo <= and_1622_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_117_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1512_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_117_sva_dfm_2_enexo <= and_1512_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_197_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1672_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_197_sva_dfm_2_enexo <= and_1672_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_71_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1420_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_71_sva_dfm_2_enexo <= and_1420_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_31_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1340_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_31_sva_dfm_2_enexo <= and_1340_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_41_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1360_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_41_sva_dfm_2_enexo <= and_1360_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_158_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1594_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_158_sva_dfm_2_enexo <= and_1594_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_58_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1394_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_58_sva_dfm_2_enexo <= and_1394_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_76_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1430_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_76_sva_dfm_2_enexo <= and_1430_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_24_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1326_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_24_sva_dfm_2_enexo <= and_1326_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_65_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1408_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_65_sva_dfm_2_enexo <= and_1408_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_40_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1358_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_40_sva_dfm_2_enexo <= and_1358_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_30_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1338_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_30_sva_dfm_2_enexo <= and_1338_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_151_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1580_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_151_sva_dfm_2_enexo <= and_1580_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_44_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1366_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_44_sva_dfm_2_enexo <= and_1366_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_107_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1492_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_107_sva_dfm_2_enexo <= and_1492_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_1_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1280_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_1_sva_dfm_2_enexo <= and_1280_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_39_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1356_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_39_sva_dfm_2_enexo <= and_1356_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_61_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1400_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_61_sva_dfm_2_enexo <= and_1400_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_137_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1552_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_137_sva_dfm_2_enexo <= and_1552_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_222_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1722_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_222_sva_dfm_2_enexo <= and_1722_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_165_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1608_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_165_sva_dfm_2_enexo <= and_1608_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_94_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1466_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_94_sva_dfm_2_enexo <= and_1466_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_254_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1786_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_254_sva_dfm_2_enexo <= and_1786_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_207_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1692_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_207_sva_dfm_2_enexo <= and_1692_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_47_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1372_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_47_sva_dfm_2_enexo <= and_1372_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_89_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1456_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_89_sva_dfm_2_enexo <= and_1456_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_228_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1734_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_228_sva_dfm_2_enexo <= and_1734_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_234_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1746_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_234_sva_dfm_2_enexo <= and_1746_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_193_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1664_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_193_sva_dfm_2_enexo <= and_1664_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_187_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1652_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_187_sva_dfm_2_enexo <= and_1652_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_45_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1368_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_45_sva_dfm_2_enexo <= and_1368_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_112_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1502_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_112_sva_dfm_2_enexo <= and_1502_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_11_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1300_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_11_sva_dfm_2_enexo <= and_1300_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_66_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1410_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_66_sva_dfm_2_enexo <= and_1410_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_15_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1308_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_15_sva_dfm_2_enexo <= and_1308_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1_enexo
          <= 1'b1;
    end
    else if ( rva_in_reg_rw_and_6_cse | input_mem_banks_read_1_read_data_and_5_enex5
        ) begin
      reg_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1_enexo
          <= rva_in_reg_rw_and_6_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_184_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1646_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_184_sva_dfm_2_enexo <= and_1646_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_103_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1484_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_103_sva_dfm_2_enexo <= and_1484_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_124_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1526_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_124_sva_dfm_2_enexo <= and_1526_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_182_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1642_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_182_sva_dfm_2_enexo <= and_1642_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_247_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1772_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_247_sva_dfm_2_enexo <= and_1772_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_84_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1446_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_84_sva_dfm_2_enexo <= and_1446_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_167_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1612_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_167_sva_dfm_2_enexo <= and_1612_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_148_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1574_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_148_sva_dfm_2_enexo <= and_1574_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_227_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1732_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_227_sva_dfm_2_enexo <= and_1732_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_232_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1742_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_232_sva_dfm_2_enexo <= and_1742_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_186_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1650_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_186_sva_dfm_2_enexo <= and_1650_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_253_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1784_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_253_sva_dfm_2_enexo <= and_1784_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_105_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1488_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_105_sva_dfm_2_enexo <= and_1488_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_101_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1480_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_101_sva_dfm_2_enexo <= and_1480_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_7_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1292_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_7_sva_dfm_2_enexo <= and_1292_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_5_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1288_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_5_sva_dfm_2_enexo <= and_1288_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_201_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1680_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_201_sva_dfm_2_enexo <= and_1680_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_236_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1750_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_236_sva_dfm_2_enexo <= and_1750_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_195_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1668_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_195_sva_dfm_2_enexo <= and_1668_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_62_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1402_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_62_sva_dfm_2_enexo <= and_1402_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_92_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1462_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_92_sva_dfm_2_enexo <= and_1462_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_18_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1314_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_18_sva_dfm_2_enexo <= and_1314_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_35_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1348_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_35_sva_dfm_2_enexo <= and_1348_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_210_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1698_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_210_sva_dfm_2_enexo <= and_1698_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_106_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1490_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_106_sva_dfm_2_enexo <= and_1490_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_70_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1418_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_70_sva_dfm_2_enexo <= and_1418_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_126_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1530_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_126_sva_dfm_2_enexo <= and_1530_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_sva_1_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_30_tmp | input_mem_banks_read_1_read_data_and_5_enex5
        ) begin
      reg_input_mem_banks_read_read_data_sva_1_enexo <= input_mem_banks_read_read_data_and_30_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_3_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1284_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_3_sva_dfm_2_enexo <= and_1284_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_97_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1472_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_97_sva_dfm_2_enexo <= and_1472_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_252_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1782_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_252_sva_dfm_2_enexo <= and_1782_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_77_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1432_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_77_sva_dfm_2_enexo <= and_1432_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_57_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1392_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_57_sva_dfm_2_enexo <= and_1392_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_217_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1712_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_217_sva_dfm_2_enexo <= and_1712_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_163_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1604_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_163_sva_dfm_2_enexo <= and_1604_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_16_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1310_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_16_sva_dfm_2_enexo <= and_1310_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_42_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1362_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_42_sva_dfm_2_enexo <= and_1362_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_219_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1716_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_219_sva_dfm_2_enexo <= and_1716_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_225_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1728_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_225_sva_dfm_2_enexo <= and_1728_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_120_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1518_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_120_sva_dfm_2_enexo <= and_1518_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_63_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1404_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_63_sva_dfm_2_enexo <= and_1404_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_229_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1736_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_229_sva_dfm_2_enexo <= and_1736_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_176_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1630_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_176_sva_dfm_2_enexo <= and_1630_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_54_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1386_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_54_sva_dfm_2_enexo <= and_1386_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_74_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1426_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_74_sva_dfm_2_enexo <= and_1426_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_80_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1438_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_80_sva_dfm_2_enexo <= and_1438_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_78_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1434_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_78_sva_dfm_2_enexo <= and_1434_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_140_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1558_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_140_sva_dfm_2_enexo <= and_1558_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_153_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1584_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_153_sva_dfm_2_enexo <= and_1584_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_174_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1626_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_174_sva_dfm_2_enexo <= and_1626_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_156_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1590_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_156_sva_dfm_2_enexo <= and_1590_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_202_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1682_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_202_sva_dfm_2_enexo <= and_1682_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_238_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1754_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_238_sva_dfm_2_enexo <= and_1754_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_67_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1412_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_67_sva_dfm_2_enexo <= and_1412_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_87_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1452_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_87_sva_dfm_2_enexo <= and_1452_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_147_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1572_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_147_sva_dfm_2_enexo <= and_1572_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_170_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1618_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_170_sva_dfm_2_enexo <= and_1618_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_2_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1282_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_2_sva_dfm_2_enexo <= and_1282_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_29_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1336_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_29_sva_dfm_2_enexo <= and_1336_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_183_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1644_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_183_sva_dfm_2_enexo <= and_1644_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_166_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1610_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_166_sva_dfm_2_enexo <= and_1610_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_33_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1344_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_33_sva_dfm_2_enexo <= and_1344_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_134_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1546_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_134_sva_dfm_2_enexo <= and_1546_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_162_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1602_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_162_sva_dfm_2_enexo <= and_1602_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_159_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1596_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_159_sva_dfm_2_enexo <= and_1596_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_51_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1380_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_51_sva_dfm_2_enexo <= and_1380_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_152_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1582_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_152_sva_dfm_2_enexo <= and_1582_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_173_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1624_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_173_sva_dfm_2_enexo <= and_1624_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_179_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1636_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_179_sva_dfm_2_enexo <= and_1636_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_180_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1638_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_180_sva_dfm_2_enexo <= and_1638_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_144_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1566_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_144_sva_dfm_2_enexo <= and_1566_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_209_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1696_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_209_sva_dfm_2_enexo <= and_1696_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_48_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1374_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_48_sva_dfm_2_enexo <= and_1374_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_160_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1598_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_160_sva_dfm_2_enexo <= and_1598_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_203_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1684_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_203_sva_dfm_2_enexo <= and_1684_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_20_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1318_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_20_sva_dfm_2_enexo <= and_1318_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_43_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1364_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_43_sva_dfm_2_enexo <= and_1364_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_237_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1752_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_237_sva_dfm_2_enexo <= and_1752_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_102_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1482_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_102_sva_dfm_2_enexo <= and_1482_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_111_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1500_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_111_sva_dfm_2_enexo <= and_1500_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_129_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1536_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_129_sva_dfm_2_enexo <= and_1536_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_100_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1478_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_100_sva_dfm_2_enexo <= and_1478_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_10_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1298_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_10_sva_dfm_2_enexo <= and_1298_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_145_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1568_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_145_sva_dfm_2_enexo <= and_1568_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_239_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1756_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_239_sva_dfm_2_enexo <= and_1756_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_196_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1670_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_196_sva_dfm_2_enexo <= and_1670_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_56_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1390_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_56_sva_dfm_2_enexo <= and_1390_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_154_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1586_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_154_sva_dfm_2_enexo <= and_1586_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_141_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1560_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_141_sva_dfm_2_enexo <= and_1560_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_245_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1768_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_245_sva_dfm_2_enexo <= and_1768_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_128_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1534_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_128_sva_dfm_2_enexo <= and_1534_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_164_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1606_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_164_sva_dfm_2_enexo <= and_1606_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_175_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1628_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_175_sva_dfm_2_enexo <= and_1628_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_69_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1416_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_69_sva_dfm_2_enexo <= and_1416_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_6_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1290_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_6_sva_dfm_2_enexo <= and_1290_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_125_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1528_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_125_sva_dfm_2_enexo <= and_1528_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_127_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1532_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_127_sva_dfm_2_enexo <= and_1532_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_82_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1442_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_82_sva_dfm_2_enexo <= and_1442_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_25_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1328_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_25_sva_dfm_2_enexo <= and_1328_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_226_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1730_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_226_sva_dfm_2_enexo <= and_1730_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_138_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1554_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_138_sva_dfm_2_enexo <= and_1554_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_133_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1544_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_133_sva_dfm_2_enexo <= and_1544_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_37_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1352_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_37_sva_dfm_2_enexo <= and_1352_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_242_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1762_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_242_sva_dfm_2_enexo <= and_1762_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_171_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1620_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_171_sva_dfm_2_enexo <= and_1620_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_216_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1710_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_216_sva_dfm_2_enexo <= and_1710_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_206_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1690_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_206_sva_dfm_2_enexo <= and_1690_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_9_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1296_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_9_sva_dfm_2_enexo <= and_1296_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_32_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1342_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_32_sva_dfm_2_enexo <= and_1342_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_86_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1450_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_86_sva_dfm_2_enexo <= and_1450_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_122_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1522_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_122_sva_dfm_2_enexo <= and_1522_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_26_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1330_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_26_sva_dfm_2_enexo <= and_1330_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_190_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1658_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_190_sva_dfm_2_enexo <= and_1658_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_199_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1676_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_199_sva_dfm_2_enexo <= and_1676_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_73_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1424_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_73_sva_dfm_2_enexo <= and_1424_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_79_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1436_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_79_sva_dfm_2_enexo <= and_1436_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_114_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1506_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_114_sva_dfm_2_enexo <= and_1506_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_131_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1540_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_131_sva_dfm_2_enexo <= and_1540_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_198_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1674_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_198_sva_dfm_2_enexo <= and_1674_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_98_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1474_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_98_sva_dfm_2_enexo <= and_1474_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_168_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1614_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_168_sva_dfm_2_enexo <= and_1614_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_146_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1570_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_146_sva_dfm_2_enexo <= and_1570_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_211_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1700_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_211_sva_dfm_2_enexo <= and_1700_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_233_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1744_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_233_sva_dfm_2_enexo <= and_1744_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_115_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1508_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_115_sva_dfm_2_enexo <= and_1508_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_215_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1708_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_215_sva_dfm_2_enexo <= and_1708_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_212_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1702_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_212_sva_dfm_2_enexo <= and_1702_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_200_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1678_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_200_sva_dfm_2_enexo <= and_1678_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_143_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1564_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_143_sva_dfm_2_enexo <= and_1564_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_185_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1648_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_185_sva_dfm_2_enexo <= and_1648_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_23_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1324_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_23_sva_dfm_2_enexo <= and_1324_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_205_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1688_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_205_sva_dfm_2_enexo <= and_1688_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_99_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1476_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_99_sva_dfm_2_enexo <= and_1476_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_38_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1354_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_38_sva_dfm_2_enexo <= and_1354_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_230_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1738_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_230_sva_dfm_2_enexo <= and_1738_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_218_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1714_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_218_sva_dfm_2_enexo <= and_1714_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_244_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1766_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_244_sva_dfm_2_enexo <= and_1766_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_161_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1600_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_161_sva_dfm_2_enexo <= and_1600_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_60_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1398_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_60_sva_dfm_2_enexo <= and_1398_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_130_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1538_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_130_sva_dfm_2_enexo <= and_1538_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_178_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1634_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_178_sva_dfm_2_enexo <= and_1634_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_119_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1516_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_119_sva_dfm_2_enexo <= and_1516_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_118_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1514_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_118_sva_dfm_2_enexo <= and_1514_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_34_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1346_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_34_sva_dfm_2_enexo <= and_1346_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_28_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1334_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_28_sva_dfm_2_enexo <= and_1334_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_85_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1448_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_85_sva_dfm_2_enexo <= and_1448_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_64_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1406_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_64_sva_dfm_2_enexo <= and_1406_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_59_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1396_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_59_sva_dfm_2_enexo <= and_1396_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_0_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1278_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_0_sva_dfm_2_enexo <= and_1278_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_50_enex5 | rva_out_reg_data_and_104_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_4_enexo <= rva_out_reg_data_and_50_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1792_cse | rva_out_reg_data_and_105_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= and_1792_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1792_cse | rva_out_reg_data_and_106_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo <= and_1792_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_29_tmp | input_mem_banks_read_read_data_and_28_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_read_data_and_29_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( weight_mem_banks_load_store_for_else_and_17_ssc | rva_out_reg_data_and_50_enex5
        ) begin
      reg_weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_1_enexo
          <= weight_mem_banks_load_store_for_else_and_17_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_70_cse | rva_out_reg_data_and_107_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= rva_out_reg_data_and_70_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_70_cse | rva_out_reg_data_and_108_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= rva_out_reg_data_and_70_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_115_enex5 | rva_out_reg_data_and_109_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= rva_out_reg_data_and_115_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_116_enex5 | rva_out_reg_data_and_110_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= rva_out_reg_data_and_116_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_117_enex5 | rva_out_reg_data_and_111_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= rva_out_reg_data_and_117_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_118_enex5 | rva_out_reg_data_and_112_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= rva_out_reg_data_and_118_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_119_enex5 | rva_out_reg_data_and_113_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo <= rva_out_reg_data_and_119_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_120_enex5 | rva_out_reg_data_and_114_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo <= rva_out_reg_data_and_120_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_78_enex5 | rva_out_reg_data_and_115_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= rva_out_reg_data_and_78_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_121_enex5 | rva_out_reg_data_and_116_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= rva_out_reg_data_and_121_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_122_enex5 | rva_out_reg_data_and_117_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= rva_out_reg_data_and_122_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_123_enex5 | rva_out_reg_data_and_118_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= rva_out_reg_data_and_123_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_124_enex5 | rva_out_reg_data_and_119_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo <= rva_out_reg_data_and_124_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_125_enex5 | rva_out_reg_data_and_120_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo <= rva_out_reg_data_and_125_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse | rva_out_reg_data_and_78_enex5
        ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_85_cse | rva_out_reg_data_and_121_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= rva_out_reg_data_and_85_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_85_cse | rva_out_reg_data_and_122_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= rva_out_reg_data_and_85_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_85_cse | rva_out_reg_data_and_123_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= rva_out_reg_data_and_85_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_85_cse | rva_out_reg_data_and_124_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo <= rva_out_reg_data_and_85_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_85_cse | rva_out_reg_data_and_125_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_1_enexo <= rva_out_reg_data_and_85_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_101_enex5 | weight_port_read_out_data_and_99_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_101_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_102_enex5 | weight_port_read_out_data_and_100_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_enexo <= weight_port_read_out_data_and_102_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_131_enex5 | rva_out_reg_data_and_126_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_1_enexo <= rva_out_reg_data_and_131_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_132_enex5 | rva_out_reg_data_and_127_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_1_enexo <= rva_out_reg_data_and_132_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_133_enex5 | rva_out_reg_data_and_128_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_133_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_134_enex5 | rva_out_reg_data_and_129_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo <= rva_out_reg_data_and_134_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_135_enex5 | rva_out_reg_data_and_130_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_135_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_94_ssc | rva_out_reg_data_and_131_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo <= weight_port_read_out_data_and_94_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_17_itm_1_2_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_222_ssc | rva_out_reg_data_and_132_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_17_itm_1_2_enexo <= weight_mem_run_3_for_5_and_222_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_ssc | weight_port_read_out_data_and_101_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_15_8_4_itm_1_1_enexo
          <= input_mem_banks_read_1_read_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_ssc | weight_port_read_out_data_and_102_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_slc_input_mem_banks_read_1_read_data_7_0_3_itm_1_1_enexo
          <= input_mem_banks_read_1_read_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( and_1792_cse | rva_out_reg_data_and_133_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_1_enexo <= and_1792_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1792_cse | rva_out_reg_data_and_134_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo <= and_1792_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( and_1792_cse | rva_out_reg_data_and_135_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_1_enexo <= and_1792_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_105_enex5 | weight_port_read_out_data_and_103_enex5
        ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo <= weight_port_read_out_data_and_105_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_106_enex5 | weight_port_read_out_data_and_104_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_2_enexo <= weight_port_read_out_data_and_106_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_17_itm_1_2_enexo_1 <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_222_ssc | weight_port_read_out_data_and_105_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_17_itm_1_2_enexo_1 <= weight_mem_run_3_for_5_and_222_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo_1 <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_94_ssc | weight_port_read_out_data_and_106_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo_1 <= weight_port_read_out_data_and_94_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_95_enex5 | rva_out_reg_data_and_136_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_9_1_enexo <= rva_out_reg_data_and_95_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_94_enex5 | rva_out_reg_data_and_137_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_7_1_enexo <= rva_out_reg_data_and_94_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_99_enex5 | rva_out_reg_data_and_138_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_enexo <= rva_out_reg_data_and_99_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_100_enex5 | rva_out_reg_data_and_139_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_1_enexo <= rva_out_reg_data_and_100_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_97_enex5 | rva_out_reg_data_and_140_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_1_enexo <= rva_out_reg_data_and_97_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_95_enex5 | weight_port_read_out_data_and_107_enex5
        ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_1_enexo
          <= weight_port_read_out_data_and_95_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_1_enexo
          <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_96_enex5 | weight_port_read_out_data_and_108_enex5
        ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_1_enexo
          <= weight_port_read_out_data_and_96_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_2_enexo
          <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_97_enex5 | weight_port_read_out_data_and_109_enex5
        ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_2_enexo
          <= weight_port_read_out_data_and_97_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_98_enex5 | weight_port_read_out_data_and_110_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_2_enexo <= weight_port_read_out_data_and_98_enex5;
    end
  end
  assign nl_operator_4_false_acc_nl = pe_config_manager_counter_sva_mx1 + 4'b0001;
  assign operator_4_false_acc_nl = nl_operator_4_false_acc_nl[3:0];
  assign pe_config_UpdateManagerCounter_if_not_7_nl = ~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  assign nl_input_read_addrs_sva_1_1  = pe_config_input_counter_sva_mx1 + pe_manager_base_input_sva_mx1_7_0;
  assign PECore_RunScale_if_for_3_scaled_val_mul_1_nl = (accum_vector_data_2_18_0_sva)
      * 8'b10100111;
  assign or_418_nl = PECore_RunMac_PECore_RunMac_if_and_svs_st_9 | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_9);
  assign nor_296_nl = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3) | rva_in_reg_rw_sva_4);
  assign mux_5_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_3_lpi_1_dfm_1, nor_296_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign nor_297_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_run_3_for_land_3_lpi_1_dfm_1));
  assign mux_6_nl = MUX_s_1_2_2(mux_5_nl, nor_297_nl, or_tmp_2);
  assign or_12_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp;
  assign mux_7_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_5_lpi_1_dfm_1, or_12_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_11_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_5_lpi_1_dfm_1;
  assign or_10_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1;
  assign mux_8_nl = MUX_s_1_2_2(mux_7_nl, or_11_nl, or_10_nl);
  assign mux_9_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_7_lpi_1_dfm_1, (~ rva_in_reg_rw_sva_4),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_run_3_for_5_and_100_nl = (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_lpi_1_dfm_1;
  assign mux_31_nl = MUX_s_1_2_2(or_tmp_60, (~ or_38_cse), rva_in_reg_rw_sva_st_1_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_20_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_76_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[7:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_76_nl);
  assign nor_nl = ~((~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_32_nl = MUX_s_1_2_2(nor_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_72_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[7:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_72_nl);
  assign nor_298_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_69_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1));
  assign mux_33_nl = MUX_s_1_2_2(nor_298_nl, or_69_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1);
  assign or_76_nl = (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])))
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign or_74_nl = (~(and_706_cse | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1))
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_34_nl = MUX_s_1_2_2(or_76_nl, or_74_nl, while_stage_0_5);
  assign or_71_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_35_nl = MUX_s_1_2_2(mux_34_nl, or_71_nl, while_stage_0_6);
  assign nor_303_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ while_stage_0_6));
  assign mux_36_nl = MUX_s_1_2_2(nor_303_nl, while_stage_0_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_78_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & while_stage_0_6));
  assign or_77_nl = (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
      | (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign mux_37_nl = MUX_s_1_2_2(mux_36_nl, or_78_nl, or_77_nl);
  assign mux_38_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_3, (weight_mem_write_arbxbar_xbar_for_empty_sva_1[3]),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign nor_700_nl = ~((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign nor_701_nl = ~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | (~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse)));
  assign mux_359_nl = MUX_s_1_2_2(nor_700_nl, nor_701_nl, while_stage_0_3);
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2,
      while_stage_0_4);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl
      = MUX_v_11_2_2(11'b00000000000, PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl
      = MUX_v_4_2_2(4'b0000, pe_config_manager_counter_sva_mx1, PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign and_600_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & and_dcpl_203 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]));
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl = (state_mux_1_cse!=2'b00)
      | state_0_sva_mx1;
  assign PECore_UpdateFSM_switch_lp_or_nl = PECore_UpdateFSM_switch_lp_equal_tmp_6
      | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  assign PECore_UpdateFSM_switch_lp_mux1h_15_nl = MUX1HOT_v_2_3_2((signext_2_1(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl)),
      2'b01, 2'b10, {PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      , PECore_UpdateFSM_switch_lp_or_nl , PECore_RunScale_PECore_RunScale_if_and_1_svs_1});
  assign PECore_UpdateFSM_switch_lp_nor_8_nl = ~(PECore_PushOutput_PECore_PushOutput_if_and_svs_1
      | PECore_UpdateFSM_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_and_1_nl = MUX_v_2_2_2(2'b00, PECore_UpdateFSM_switch_lp_mux1h_15_nl,
      PECore_UpdateFSM_switch_lp_nor_8_nl);
  assign nor_712_nl = ~((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | (~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1);
  assign nand_241_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & ((~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1));
  assign mux_361_nl = MUX_s_1_2_2(nor_712_nl, nand_241_nl, PECore_UpdateFSM_switch_lp_equal_tmp_3_1);
  assign nor_713_nl = ~((~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1);
  assign mux_362_nl = MUX_s_1_2_2(and_1884_cse, nor_713_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nl_operator_8_false_acc_sdt_sva_1  = conv_u2s_8_9(pe_config_num_output_sva)
      + 9'b111111111;
  assign nl_ProductSum_for_acc_23_nl = conv_u2u_18_19(Datapath_for_3_ProductSum_for_acc_3_1)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_21_z);
  assign ProductSum_for_acc_23_nl = nl_ProductSum_for_acc_23_nl[18:0];
  assign nl_ProductSum_for_acc_21_nl = ProductSum_for_acc_22_itm_1 + ProductSum_for_acc_23_nl;
  assign ProductSum_for_acc_21_nl = nl_ProductSum_for_acc_21_nl[18:0];
  assign PECore_UpdateFSM_switch_lp_not_19_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_129_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_115_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_122_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_94_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_108_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_130_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_131_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_133_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign and_922_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])
      & (~ or_713_tmp);
  assign and_923_nl = and_dcpl_596 & (~ or_713_tmp);
  assign and_924_nl = nor_260_cse & (~ or_713_tmp);
  assign mux1h_1_nl = MUX1HOT_v_8_3_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[63:56]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[63:56]), (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[15:8]),
      {and_922_nl , and_923_nl , and_924_nl});
  assign not_2217_nl = ~ or_713_tmp;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_123_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_126_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_127_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_128_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_109_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_110_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_112_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_114_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign and_610_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign and_612_nl = and_dcpl_599 & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign and_616_nl = and_dcpl_603 & (~(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4));
  assign and_620_nl = (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      & weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_621_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_load_store_for_else_mux1h_17_nl = MUX1HOT_v_8_5_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[47:40]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[47:40]), (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[7:0]),
      (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[7:0]), (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[7:0]),
      {and_610_nl , and_612_nl , and_616_nl , and_620_nl , and_621_nl});
  assign and_613_nl = and_dcpl_599 & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]));
  assign weight_mem_banks_load_store_for_else_or_nl = MUX_v_8_2_2(weight_mem_banks_load_store_for_else_mux1h_17_nl,
      8'b11111111, and_613_nl);
  assign or_715_nl = ((~((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]) | (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2])))
      & and_dcpl_599) | ((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & and_dcpl_603 & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_321_nl = MUX_v_8_2_2(weight_mem_banks_load_store_for_else_or_nl, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[7:0]),
      or_715_nl);
  assign mux_307_nl = MUX_s_1_2_2((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]),
      (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign nor_425_nl = ~((mux_307_nl & and_dcpl_599) | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[2])
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])));
  assign mux_65_nl = MUX_s_1_2_2(or_tmp_94, (~ or_tmp_95), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign mux_64_nl = MUX_s_1_2_2((~ or_tmp_95), or_tmp_94, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign mux_66_nl = MUX_s_1_2_2(mux_65_nl, mux_64_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_63_nl = MUX_s_1_2_2((~ or_tmp_95), or_tmp_94, or_231_cse);
  assign mux_67_nl = MUX_s_1_2_2(mux_66_nl, mux_63_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_68_nl = MUX_s_1_2_2(or_tmp_94, mux_67_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_124_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_125_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_132_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_78_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_111_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_113_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign or_244_nl = (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse);
  assign and_236_nl = while_stage_0_5 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse));
  assign nor_31_nl = ~((~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_23_tmp));
  assign mux_71_nl = MUX_s_1_2_2(or_244_nl, and_236_nl, nor_31_nl);
  assign nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_13_nl
      = MUX_s_1_2_2(nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_5_mux_2_mx0w3,
      nvhls_leading_ones_4U_nvhls_nvhls_t_4U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_4_mux_2_mx0w2,
      operator_4_false_2_operator_4_false_2_or_mdf_3_sva_1);
  assign nand_36_nl = ~(nvhls_leading_ones_8U_nvhls_nvhls_t_8U_nvuint_t_nvhls_nvhls_t_3U_nvuint_t_1_mux_13_nl
      & operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1);
  assign or_248_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse);
  assign mux_72_nl = MUX_s_1_2_2(nand_36_nl, or_248_nl, while_stage_0_5);
  assign or_247_nl = (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse);
  assign or_245_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_operator_7_false_1_operator_7_false_1_or_tmp
      | (~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign mux_73_nl = MUX_s_1_2_2(mux_72_nl, or_247_nl, or_245_nl);
  assign or_251_nl = (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse);
  assign and_238_nl = while_stage_0_5 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse));
  assign nor_32_nl = ~((~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_7_tmp));
  assign mux_74_nl = MUX_s_1_2_2(or_251_nl, and_238_nl, nor_32_nl);
  assign or_254_nl = (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse);
  assign and_239_nl = while_stage_0_5 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_cse));
  assign nor_33_nl = ~((~ while_stage_0_4) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_3_tmp));
  assign mux_75_nl = MUX_s_1_2_2(or_254_nl, and_239_nl, nor_33_nl);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl
      = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]), pe_config_is_zero_first_sva_mx1,
      PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_19_nl
      = MUX_s_1_2_2(PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl,
      pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_or_5_cse_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b110)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b011)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b101)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_nl = (pe_manager_base_weight_sva[1])
      & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 & (~ (pe_manager_base_weight_sva[2]))
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1
      & (pe_manager_base_weight_sva[0]) & (~ (pe_manager_base_weight_sva[2])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign mux_76_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, (~ rva_in_reg_rw_sva_st_1_3),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign PECore_RunScale_if_for_1_scaled_val_mul_1_nl = (accum_vector_data_0_18_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_2_scaled_val_mul_1_nl = (accum_vector_data_1_18_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_4_scaled_val_mul_1_nl = (accum_vector_data_3_18_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_5_scaled_val_mul_1_nl = (accum_vector_data_4_18_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_6_scaled_val_mul_1_nl = (accum_vector_data_5_18_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_7_scaled_val_mul_1_nl = (accum_vector_data_6_18_0_sva)
      * 8'b10100111;
  assign PECore_RunScale_if_for_8_scaled_val_mul_1_nl = (accum_vector_data_7_18_0_sva)
      * 8'b10100111;
  assign nor_307_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | weight_mem_run_3_for_weight_mem_run_3_for_and_4_cse);
  assign mux_77_nl = MUX_s_1_2_2(or_tmp_111, nor_307_nl, weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1);
  assign mux_78_nl = MUX_s_1_2_2(mux_77_nl, or_tmp_111, weight_mem_write_arbxbar_xbar_for_empty_sva_1[6]);
  assign nl_ProductSum_for_acc_22_itm_1  = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_24_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_23_z);
  assign nl_ProductSum_for_acc_36_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_4_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_3_z);
  assign ProductSum_for_acc_36_nl = nl_ProductSum_for_acc_36_nl[18:0];
  assign nl_ProductSum_for_acc_37_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_2_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_1_z);
  assign ProductSum_for_acc_37_nl = nl_ProductSum_for_acc_37_nl[18:0];
  assign nl_ProductSum_for_acc_nl = ProductSum_for_acc_36_nl + ProductSum_for_acc_37_nl;
  assign ProductSum_for_acc_nl = nl_ProductSum_for_acc_nl[18:0];
  assign PECore_UpdateFSM_switch_lp_not_32_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign nl_ProductSum_for_acc_34_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_8_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_7_z);
  assign ProductSum_for_acc_34_nl = nl_ProductSum_for_acc_34_nl[18:0];
  assign nl_ProductSum_for_acc_35_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_6_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_5_z);
  assign ProductSum_for_acc_35_nl = nl_ProductSum_for_acc_35_nl[18:0];
  assign nl_ProductSum_for_acc_33_nl = ProductSum_for_acc_34_nl + ProductSum_for_acc_35_nl;
  assign ProductSum_for_acc_33_nl = nl_ProductSum_for_acc_33_nl[18:0];
  assign PECore_UpdateFSM_switch_lp_not_21_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign nl_ProductSum_for_acc_31_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_12_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_11_z);
  assign ProductSum_for_acc_31_nl = nl_ProductSum_for_acc_31_nl[18:0];
  assign nl_ProductSum_for_acc_32_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_10_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_9_z);
  assign ProductSum_for_acc_32_nl = nl_ProductSum_for_acc_32_nl[18:0];
  assign nl_ProductSum_for_acc_30_nl = ProductSum_for_acc_31_nl + ProductSum_for_acc_32_nl;
  assign ProductSum_for_acc_30_nl = nl_ProductSum_for_acc_30_nl[18:0];
  assign PECore_UpdateFSM_switch_lp_not_33_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign nl_ProductSum_for_acc_28_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_16_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_15_z);
  assign ProductSum_for_acc_28_nl = nl_ProductSum_for_acc_28_nl[18:0];
  assign nl_ProductSum_for_acc_29_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_14_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_13_z);
  assign ProductSum_for_acc_29_nl = nl_ProductSum_for_acc_29_nl[18:0];
  assign nl_ProductSum_for_acc_27_nl = ProductSum_for_acc_28_nl + ProductSum_for_acc_29_nl;
  assign ProductSum_for_acc_27_nl = nl_ProductSum_for_acc_27_nl[18:0];
  assign PECore_UpdateFSM_switch_lp_not_37_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign nl_ProductSum_for_acc_25_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_20_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_19_z);
  assign ProductSum_for_acc_25_nl = nl_ProductSum_for_acc_25_nl[18:0];
  assign nl_ProductSum_for_acc_26_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_18_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_17_z);
  assign ProductSum_for_acc_26_nl = nl_ProductSum_for_acc_26_nl[18:0];
  assign nl_ProductSum_for_acc_24_nl = ProductSum_for_acc_25_nl + ProductSum_for_acc_26_nl;
  assign ProductSum_for_acc_24_nl = nl_ProductSum_for_acc_24_nl[18:0];
  assign PECore_UpdateFSM_switch_lp_not_34_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign nl_ProductSum_for_acc_19_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_28_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_27_z);
  assign ProductSum_for_acc_19_nl = nl_ProductSum_for_acc_19_nl[18:0];
  assign nl_ProductSum_for_acc_20_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_26_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_25_z);
  assign ProductSum_for_acc_20_nl = nl_ProductSum_for_acc_20_nl[18:0];
  assign nl_ProductSum_for_acc_18_nl = ProductSum_for_acc_19_nl + ProductSum_for_acc_20_nl;
  assign ProductSum_for_acc_18_nl = nl_ProductSum_for_acc_18_nl[18:0];
  assign PECore_UpdateFSM_switch_lp_not_35_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign nl_ProductSum_for_acc_16_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_31_z);
  assign ProductSum_for_acc_16_nl = nl_ProductSum_for_acc_16_nl[18:0];
  assign nl_ProductSum_for_acc_17_nl = conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_30_z)
      + conv_u2u_18_19(Datapath_for_4_ProductSum_for_acc_5_cmp_29_z);
  assign ProductSum_for_acc_17_nl = nl_ProductSum_for_acc_17_nl[18:0];
  assign nl_ProductSum_for_acc_15_nl = ProductSum_for_acc_16_nl + ProductSum_for_acc_17_nl;
  assign ProductSum_for_acc_15_nl = nl_ProductSum_for_acc_15_nl[18:0];
  assign PECore_UpdateFSM_switch_lp_not_36_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  assign input_mem_banks_read_1_for_mux_4_nl = MUX_v_64_256_2(input_mem_banks_bank_a_0_sva_dfm_2,
      input_mem_banks_bank_a_1_sva_dfm_2, input_mem_banks_bank_a_2_sva_dfm_2, input_mem_banks_bank_a_3_sva_dfm_2,
      input_mem_banks_bank_a_4_sva_dfm_2, input_mem_banks_bank_a_5_sva_dfm_2, input_mem_banks_bank_a_6_sva_dfm_2,
      input_mem_banks_bank_a_7_sva_dfm_2, input_mem_banks_bank_a_8_sva_dfm_2, input_mem_banks_bank_a_9_sva_dfm_2,
      input_mem_banks_bank_a_10_sva_dfm_2, input_mem_banks_bank_a_11_sva_dfm_2, input_mem_banks_bank_a_12_sva_dfm_2,
      input_mem_banks_bank_a_13_sva_dfm_2, input_mem_banks_bank_a_14_sva_dfm_2, input_mem_banks_bank_a_15_sva_dfm_2,
      input_mem_banks_bank_a_16_sva_dfm_2, input_mem_banks_bank_a_17_sva_dfm_2, input_mem_banks_bank_a_18_sva_dfm_2,
      input_mem_banks_bank_a_19_sva_dfm_2, input_mem_banks_bank_a_20_sva_dfm_2, input_mem_banks_bank_a_21_sva_dfm_2,
      input_mem_banks_bank_a_22_sva_dfm_2, input_mem_banks_bank_a_23_sva_dfm_2, input_mem_banks_bank_a_24_sva_dfm_2,
      input_mem_banks_bank_a_25_sva_dfm_2, input_mem_banks_bank_a_26_sva_dfm_2, input_mem_banks_bank_a_27_sva_dfm_2,
      input_mem_banks_bank_a_28_sva_dfm_2, input_mem_banks_bank_a_29_sva_dfm_2, input_mem_banks_bank_a_30_sva_dfm_2,
      input_mem_banks_bank_a_31_sva_dfm_2, input_mem_banks_bank_a_32_sva_dfm_2, input_mem_banks_bank_a_33_sva_dfm_2,
      input_mem_banks_bank_a_34_sva_dfm_2, input_mem_banks_bank_a_35_sva_dfm_2, input_mem_banks_bank_a_36_sva_dfm_2,
      input_mem_banks_bank_a_37_sva_dfm_2, input_mem_banks_bank_a_38_sva_dfm_2, input_mem_banks_bank_a_39_sva_dfm_2,
      input_mem_banks_bank_a_40_sva_dfm_2, input_mem_banks_bank_a_41_sva_dfm_2, input_mem_banks_bank_a_42_sva_dfm_2,
      input_mem_banks_bank_a_43_sva_dfm_2, input_mem_banks_bank_a_44_sva_dfm_2, input_mem_banks_bank_a_45_sva_dfm_2,
      input_mem_banks_bank_a_46_sva_dfm_2, input_mem_banks_bank_a_47_sva_dfm_2, input_mem_banks_bank_a_48_sva_dfm_2,
      input_mem_banks_bank_a_49_sva_dfm_2, input_mem_banks_bank_a_50_sva_dfm_2, input_mem_banks_bank_a_51_sva_dfm_2,
      input_mem_banks_bank_a_52_sva_dfm_2, input_mem_banks_bank_a_53_sva_dfm_2, input_mem_banks_bank_a_54_sva_dfm_2,
      input_mem_banks_bank_a_55_sva_dfm_2, input_mem_banks_bank_a_56_sva_dfm_2, input_mem_banks_bank_a_57_sva_dfm_2,
      input_mem_banks_bank_a_58_sva_dfm_2, input_mem_banks_bank_a_59_sva_dfm_2, input_mem_banks_bank_a_60_sva_dfm_2,
      input_mem_banks_bank_a_61_sva_dfm_2, input_mem_banks_bank_a_62_sva_dfm_2, input_mem_banks_bank_a_63_sva_dfm_2,
      input_mem_banks_bank_a_64_sva_dfm_2, input_mem_banks_bank_a_65_sva_dfm_2, input_mem_banks_bank_a_66_sva_dfm_2,
      input_mem_banks_bank_a_67_sva_dfm_2, input_mem_banks_bank_a_68_sva_dfm_2, input_mem_banks_bank_a_69_sva_dfm_2,
      input_mem_banks_bank_a_70_sva_dfm_2, input_mem_banks_bank_a_71_sva_dfm_2, input_mem_banks_bank_a_72_sva_dfm_2,
      input_mem_banks_bank_a_73_sva_dfm_2, input_mem_banks_bank_a_74_sva_dfm_2, input_mem_banks_bank_a_75_sva_dfm_2,
      input_mem_banks_bank_a_76_sva_dfm_2, input_mem_banks_bank_a_77_sva_dfm_2, input_mem_banks_bank_a_78_sva_dfm_2,
      input_mem_banks_bank_a_79_sva_dfm_2, input_mem_banks_bank_a_80_sva_dfm_2, input_mem_banks_bank_a_81_sva_dfm_2,
      input_mem_banks_bank_a_82_sva_dfm_2, input_mem_banks_bank_a_83_sva_dfm_2, input_mem_banks_bank_a_84_sva_dfm_2,
      input_mem_banks_bank_a_85_sva_dfm_2, input_mem_banks_bank_a_86_sva_dfm_2, input_mem_banks_bank_a_87_sva_dfm_2,
      input_mem_banks_bank_a_88_sva_dfm_2, input_mem_banks_bank_a_89_sva_dfm_2, input_mem_banks_bank_a_90_sva_dfm_2,
      input_mem_banks_bank_a_91_sva_dfm_2, input_mem_banks_bank_a_92_sva_dfm_2, input_mem_banks_bank_a_93_sva_dfm_2,
      input_mem_banks_bank_a_94_sva_dfm_2, input_mem_banks_bank_a_95_sva_dfm_2, input_mem_banks_bank_a_96_sva_dfm_2,
      input_mem_banks_bank_a_97_sva_dfm_2, input_mem_banks_bank_a_98_sva_dfm_2, input_mem_banks_bank_a_99_sva_dfm_2,
      input_mem_banks_bank_a_100_sva_dfm_2, input_mem_banks_bank_a_101_sva_dfm_2,
      input_mem_banks_bank_a_102_sva_dfm_2, input_mem_banks_bank_a_103_sva_dfm_2,
      input_mem_banks_bank_a_104_sva_dfm_2, input_mem_banks_bank_a_105_sva_dfm_2,
      input_mem_banks_bank_a_106_sva_dfm_2, input_mem_banks_bank_a_107_sva_dfm_2,
      input_mem_banks_bank_a_108_sva_dfm_2, input_mem_banks_bank_a_109_sva_dfm_2,
      input_mem_banks_bank_a_110_sva_dfm_2, input_mem_banks_bank_a_111_sva_dfm_2,
      input_mem_banks_bank_a_112_sva_dfm_2, input_mem_banks_bank_a_113_sva_dfm_2,
      input_mem_banks_bank_a_114_sva_dfm_2, input_mem_banks_bank_a_115_sva_dfm_2,
      input_mem_banks_bank_a_116_sva_dfm_2, input_mem_banks_bank_a_117_sva_dfm_2,
      input_mem_banks_bank_a_118_sva_dfm_2, input_mem_banks_bank_a_119_sva_dfm_2,
      input_mem_banks_bank_a_120_sva_dfm_2, input_mem_banks_bank_a_121_sva_dfm_2,
      input_mem_banks_bank_a_122_sva_dfm_2, input_mem_banks_bank_a_123_sva_dfm_2,
      input_mem_banks_bank_a_124_sva_dfm_2, input_mem_banks_bank_a_125_sva_dfm_2,
      input_mem_banks_bank_a_126_sva_dfm_2, input_mem_banks_bank_a_127_sva_dfm_2,
      input_mem_banks_bank_a_128_sva_dfm_2, input_mem_banks_bank_a_129_sva_dfm_2,
      input_mem_banks_bank_a_130_sva_dfm_2, input_mem_banks_bank_a_131_sva_dfm_2,
      input_mem_banks_bank_a_132_sva_dfm_2, input_mem_banks_bank_a_133_sva_dfm_2,
      input_mem_banks_bank_a_134_sva_dfm_2, input_mem_banks_bank_a_135_sva_dfm_2,
      input_mem_banks_bank_a_136_sva_dfm_2, input_mem_banks_bank_a_137_sva_dfm_2,
      input_mem_banks_bank_a_138_sva_dfm_2, input_mem_banks_bank_a_139_sva_dfm_2,
      input_mem_banks_bank_a_140_sva_dfm_2, input_mem_banks_bank_a_141_sva_dfm_2,
      input_mem_banks_bank_a_142_sva_dfm_2, input_mem_banks_bank_a_143_sva_dfm_2,
      input_mem_banks_bank_a_144_sva_dfm_2, input_mem_banks_bank_a_145_sva_dfm_2,
      input_mem_banks_bank_a_146_sva_dfm_2, input_mem_banks_bank_a_147_sva_dfm_2,
      input_mem_banks_bank_a_148_sva_dfm_2, input_mem_banks_bank_a_149_sva_dfm_2,
      input_mem_banks_bank_a_150_sva_dfm_2, input_mem_banks_bank_a_151_sva_dfm_2,
      input_mem_banks_bank_a_152_sva_dfm_2, input_mem_banks_bank_a_153_sva_dfm_2,
      input_mem_banks_bank_a_154_sva_dfm_2, input_mem_banks_bank_a_155_sva_dfm_2,
      input_mem_banks_bank_a_156_sva_dfm_2, input_mem_banks_bank_a_157_sva_dfm_2,
      input_mem_banks_bank_a_158_sva_dfm_2, input_mem_banks_bank_a_159_sva_dfm_2,
      input_mem_banks_bank_a_160_sva_dfm_2, input_mem_banks_bank_a_161_sva_dfm_2,
      input_mem_banks_bank_a_162_sva_dfm_2, input_mem_banks_bank_a_163_sva_dfm_2,
      input_mem_banks_bank_a_164_sva_dfm_2, input_mem_banks_bank_a_165_sva_dfm_2,
      input_mem_banks_bank_a_166_sva_dfm_2, input_mem_banks_bank_a_167_sva_dfm_2,
      input_mem_banks_bank_a_168_sva_dfm_2, input_mem_banks_bank_a_169_sva_dfm_2,
      input_mem_banks_bank_a_170_sva_dfm_2, input_mem_banks_bank_a_171_sva_dfm_2,
      input_mem_banks_bank_a_172_sva_dfm_2, input_mem_banks_bank_a_173_sva_dfm_2,
      input_mem_banks_bank_a_174_sva_dfm_2, input_mem_banks_bank_a_175_sva_dfm_2,
      input_mem_banks_bank_a_176_sva_dfm_2, input_mem_banks_bank_a_177_sva_dfm_2,
      input_mem_banks_bank_a_178_sva_dfm_2, input_mem_banks_bank_a_179_sva_dfm_2,
      input_mem_banks_bank_a_180_sva_dfm_2, input_mem_banks_bank_a_181_sva_dfm_2,
      input_mem_banks_bank_a_182_sva_dfm_2, input_mem_banks_bank_a_183_sva_dfm_2,
      input_mem_banks_bank_a_184_sva_dfm_2, input_mem_banks_bank_a_185_sva_dfm_2,
      input_mem_banks_bank_a_186_sva_dfm_2, input_mem_banks_bank_a_187_sva_dfm_2,
      input_mem_banks_bank_a_188_sva_dfm_2, input_mem_banks_bank_a_189_sva_dfm_2,
      input_mem_banks_bank_a_190_sva_dfm_2, input_mem_banks_bank_a_191_sva_dfm_2,
      input_mem_banks_bank_a_192_sva_dfm_2, input_mem_banks_bank_a_193_sva_dfm_2,
      input_mem_banks_bank_a_194_sva_dfm_2, input_mem_banks_bank_a_195_sva_dfm_2,
      input_mem_banks_bank_a_196_sva_dfm_2, input_mem_banks_bank_a_197_sva_dfm_2,
      input_mem_banks_bank_a_198_sva_dfm_2, input_mem_banks_bank_a_199_sva_dfm_2,
      input_mem_banks_bank_a_200_sva_dfm_2, input_mem_banks_bank_a_201_sva_dfm_2,
      input_mem_banks_bank_a_202_sva_dfm_2, input_mem_banks_bank_a_203_sva_dfm_2,
      input_mem_banks_bank_a_204_sva_dfm_2, input_mem_banks_bank_a_205_sva_dfm_2,
      input_mem_banks_bank_a_206_sva_dfm_2, input_mem_banks_bank_a_207_sva_dfm_2,
      input_mem_banks_bank_a_208_sva_dfm_2, input_mem_banks_bank_a_209_sva_dfm_2,
      input_mem_banks_bank_a_210_sva_dfm_2, input_mem_banks_bank_a_211_sva_dfm_2,
      input_mem_banks_bank_a_212_sva_dfm_2, input_mem_banks_bank_a_213_sva_dfm_2,
      input_mem_banks_bank_a_214_sva_dfm_2, input_mem_banks_bank_a_215_sva_dfm_2,
      input_mem_banks_bank_a_216_sva_dfm_2, input_mem_banks_bank_a_217_sva_dfm_2,
      input_mem_banks_bank_a_218_sva_dfm_2, input_mem_banks_bank_a_219_sva_dfm_2,
      input_mem_banks_bank_a_220_sva_dfm_2, input_mem_banks_bank_a_221_sva_dfm_2,
      input_mem_banks_bank_a_222_sva_dfm_2, input_mem_banks_bank_a_223_sva_dfm_2,
      input_mem_banks_bank_a_224_sva_dfm_2, input_mem_banks_bank_a_225_sva_dfm_2,
      input_mem_banks_bank_a_226_sva_dfm_2, input_mem_banks_bank_a_227_sva_dfm_2,
      input_mem_banks_bank_a_228_sva_dfm_2, input_mem_banks_bank_a_229_sva_dfm_2,
      input_mem_banks_bank_a_230_sva_dfm_2, input_mem_banks_bank_a_231_sva_dfm_2,
      input_mem_banks_bank_a_232_sva_dfm_2, input_mem_banks_bank_a_233_sva_dfm_2,
      input_mem_banks_bank_a_234_sva_dfm_2, input_mem_banks_bank_a_235_sva_dfm_2,
      input_mem_banks_bank_a_236_sva_dfm_2, input_mem_banks_bank_a_237_sva_dfm_2,
      input_mem_banks_bank_a_238_sva_dfm_2, input_mem_banks_bank_a_239_sva_dfm_2,
      input_mem_banks_bank_a_240_sva_dfm_2, input_mem_banks_bank_a_241_sva_dfm_2,
      input_mem_banks_bank_a_242_sva_dfm_2, input_mem_banks_bank_a_243_sva_dfm_2,
      input_mem_banks_bank_a_244_sva_dfm_2, input_mem_banks_bank_a_245_sva_dfm_2,
      input_mem_banks_bank_a_246_sva_dfm_2, input_mem_banks_bank_a_247_sva_dfm_2,
      input_mem_banks_bank_a_248_sva_dfm_2, input_mem_banks_bank_a_249_sva_dfm_2,
      input_mem_banks_bank_a_250_sva_dfm_2, input_mem_banks_bank_a_251_sva_dfm_2,
      input_mem_banks_bank_a_252_sva_dfm_2, input_mem_banks_bank_a_253_sva_dfm_2,
      input_mem_banks_bank_a_254_sva_dfm_2, input_mem_banks_bank_a_255_sva_dfm_2,
      input_read_addrs_sva_1_1);
  assign and_633_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign weight_port_read_out_data_mux_71_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_13_mx0w2,
      weight_port_read_out_data_0_7_sva_dfm_3_7, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_135_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[15:8]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_135_nl);
  assign and_639_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign nor_418_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign while_if_while_if_and_2_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:0])
      & ({{14{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & ({{14{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
  assign or_492_nl = or_dcpl_141 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) |
      (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | or_dcpl_275;
  assign mux_90_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign mux_93_nl = MUX_s_1_2_2(nand_39_cse, rva_in_reg_rw_sva_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_404_nl = PECore_RunFSM_switch_lp_equal_tmp_1_2 & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_40_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp);
  assign or_323_nl = and_715_cse | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp;
  assign mux_94_nl = MUX_s_1_2_2(and_404_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      or_323_nl);
  assign nor_314_nl = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2) | rva_in_reg_rw_sva_3
      | input_read_req_valid_lpi_1_dfm_1_3 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1
      | rva_in_reg_rw_sva_st_1_3);
  assign mux_95_nl = MUX_s_1_2_2(mux_94_nl, nor_314_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1
      & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_1_itm_1
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2,
      (pe_manager_base_weight_sva_mx1_3_0[0]), PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_4_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2,
      (pe_manager_base_weight_sva_mx2[8]), PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl =
      (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_5_nl = MUX_s_1_2_2(pe_config_is_valid_sva,
      pe_manager_zero_active_sva, and_301_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_6_nl = MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1,
      (pe_manager_num_input_sva[0]), and_301_cse);
  assign input_mem_banks_bank_a_mux_1_nl = MUX_v_64_2_2(input_mem_banks_bank_a_0_sva_dfm_2,
      input_mem_banks_bank_a_0_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_3_nl = MUX_v_64_2_2(input_mem_banks_bank_a_1_sva_dfm_2,
      input_mem_banks_bank_a_1_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_5_nl = MUX_v_64_2_2(input_mem_banks_bank_a_2_sva_dfm_2,
      input_mem_banks_bank_a_2_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_7_nl = MUX_v_64_2_2(input_mem_banks_bank_a_3_sva_dfm_2,
      input_mem_banks_bank_a_3_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_9_nl = MUX_v_64_2_2(input_mem_banks_bank_a_4_sva_dfm_2,
      input_mem_banks_bank_a_4_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_11_nl = MUX_v_64_2_2(input_mem_banks_bank_a_5_sva_dfm_2,
      input_mem_banks_bank_a_5_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_13_nl = MUX_v_64_2_2(input_mem_banks_bank_a_6_sva_dfm_2,
      input_mem_banks_bank_a_6_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_15_nl = MUX_v_64_2_2(input_mem_banks_bank_a_7_sva_dfm_2,
      input_mem_banks_bank_a_7_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_17_nl = MUX_v_64_2_2(input_mem_banks_bank_a_8_sva_dfm_2,
      input_mem_banks_bank_a_8_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_19_nl = MUX_v_64_2_2(input_mem_banks_bank_a_9_sva_dfm_2,
      input_mem_banks_bank_a_9_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_21_nl = MUX_v_64_2_2(input_mem_banks_bank_a_10_sva_dfm_2,
      input_mem_banks_bank_a_10_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_23_nl = MUX_v_64_2_2(input_mem_banks_bank_a_11_sva_dfm_2,
      input_mem_banks_bank_a_11_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_25_nl = MUX_v_64_2_2(input_mem_banks_bank_a_12_sva_dfm_2,
      input_mem_banks_bank_a_12_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_27_nl = MUX_v_64_2_2(input_mem_banks_bank_a_13_sva_dfm_2,
      input_mem_banks_bank_a_13_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_29_nl = MUX_v_64_2_2(input_mem_banks_bank_a_14_sva_dfm_2,
      input_mem_banks_bank_a_14_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_31_nl = MUX_v_64_2_2(input_mem_banks_bank_a_15_sva_dfm_2,
      input_mem_banks_bank_a_15_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_33_nl = MUX_v_64_2_2(input_mem_banks_bank_a_16_sva_dfm_2,
      input_mem_banks_bank_a_16_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_35_nl = MUX_v_64_2_2(input_mem_banks_bank_a_17_sva_dfm_2,
      input_mem_banks_bank_a_17_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_37_nl = MUX_v_64_2_2(input_mem_banks_bank_a_18_sva_dfm_2,
      input_mem_banks_bank_a_18_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_39_nl = MUX_v_64_2_2(input_mem_banks_bank_a_19_sva_dfm_2,
      input_mem_banks_bank_a_19_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_41_nl = MUX_v_64_2_2(input_mem_banks_bank_a_20_sva_dfm_2,
      input_mem_banks_bank_a_20_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_43_nl = MUX_v_64_2_2(input_mem_banks_bank_a_21_sva_dfm_2,
      input_mem_banks_bank_a_21_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_45_nl = MUX_v_64_2_2(input_mem_banks_bank_a_22_sva_dfm_2,
      input_mem_banks_bank_a_22_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_47_nl = MUX_v_64_2_2(input_mem_banks_bank_a_23_sva_dfm_2,
      input_mem_banks_bank_a_23_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_49_nl = MUX_v_64_2_2(input_mem_banks_bank_a_24_sva_dfm_2,
      input_mem_banks_bank_a_24_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_51_nl = MUX_v_64_2_2(input_mem_banks_bank_a_25_sva_dfm_2,
      input_mem_banks_bank_a_25_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_53_nl = MUX_v_64_2_2(input_mem_banks_bank_a_26_sva_dfm_2,
      input_mem_banks_bank_a_26_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_55_nl = MUX_v_64_2_2(input_mem_banks_bank_a_27_sva_dfm_2,
      input_mem_banks_bank_a_27_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_57_nl = MUX_v_64_2_2(input_mem_banks_bank_a_28_sva_dfm_2,
      input_mem_banks_bank_a_28_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_59_nl = MUX_v_64_2_2(input_mem_banks_bank_a_29_sva_dfm_2,
      input_mem_banks_bank_a_29_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_61_nl = MUX_v_64_2_2(input_mem_banks_bank_a_30_sva_dfm_2,
      input_mem_banks_bank_a_30_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_63_nl = MUX_v_64_2_2(input_mem_banks_bank_a_31_sva_dfm_2,
      input_mem_banks_bank_a_31_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_65_nl = MUX_v_64_2_2(input_mem_banks_bank_a_32_sva_dfm_2,
      input_mem_banks_bank_a_32_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_67_nl = MUX_v_64_2_2(input_mem_banks_bank_a_33_sva_dfm_2,
      input_mem_banks_bank_a_33_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_69_nl = MUX_v_64_2_2(input_mem_banks_bank_a_34_sva_dfm_2,
      input_mem_banks_bank_a_34_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_71_nl = MUX_v_64_2_2(input_mem_banks_bank_a_35_sva_dfm_2,
      input_mem_banks_bank_a_35_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_73_nl = MUX_v_64_2_2(input_mem_banks_bank_a_36_sva_dfm_2,
      input_mem_banks_bank_a_36_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_75_nl = MUX_v_64_2_2(input_mem_banks_bank_a_37_sva_dfm_2,
      input_mem_banks_bank_a_37_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_77_nl = MUX_v_64_2_2(input_mem_banks_bank_a_38_sva_dfm_2,
      input_mem_banks_bank_a_38_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_79_nl = MUX_v_64_2_2(input_mem_banks_bank_a_39_sva_dfm_2,
      input_mem_banks_bank_a_39_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_81_nl = MUX_v_64_2_2(input_mem_banks_bank_a_40_sva_dfm_2,
      input_mem_banks_bank_a_40_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_83_nl = MUX_v_64_2_2(input_mem_banks_bank_a_41_sva_dfm_2,
      input_mem_banks_bank_a_41_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_85_nl = MUX_v_64_2_2(input_mem_banks_bank_a_42_sva_dfm_2,
      input_mem_banks_bank_a_42_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_87_nl = MUX_v_64_2_2(input_mem_banks_bank_a_43_sva_dfm_2,
      input_mem_banks_bank_a_43_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_89_nl = MUX_v_64_2_2(input_mem_banks_bank_a_44_sva_dfm_2,
      input_mem_banks_bank_a_44_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_91_nl = MUX_v_64_2_2(input_mem_banks_bank_a_45_sva_dfm_2,
      input_mem_banks_bank_a_45_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_93_nl = MUX_v_64_2_2(input_mem_banks_bank_a_46_sva_dfm_2,
      input_mem_banks_bank_a_46_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_95_nl = MUX_v_64_2_2(input_mem_banks_bank_a_47_sva_dfm_2,
      input_mem_banks_bank_a_47_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_97_nl = MUX_v_64_2_2(input_mem_banks_bank_a_48_sva_dfm_2,
      input_mem_banks_bank_a_48_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_99_nl = MUX_v_64_2_2(input_mem_banks_bank_a_49_sva_dfm_2,
      input_mem_banks_bank_a_49_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_101_nl = MUX_v_64_2_2(input_mem_banks_bank_a_50_sva_dfm_2,
      input_mem_banks_bank_a_50_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_103_nl = MUX_v_64_2_2(input_mem_banks_bank_a_51_sva_dfm_2,
      input_mem_banks_bank_a_51_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_105_nl = MUX_v_64_2_2(input_mem_banks_bank_a_52_sva_dfm_2,
      input_mem_banks_bank_a_52_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_107_nl = MUX_v_64_2_2(input_mem_banks_bank_a_53_sva_dfm_2,
      input_mem_banks_bank_a_53_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_109_nl = MUX_v_64_2_2(input_mem_banks_bank_a_54_sva_dfm_2,
      input_mem_banks_bank_a_54_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_111_nl = MUX_v_64_2_2(input_mem_banks_bank_a_55_sva_dfm_2,
      input_mem_banks_bank_a_55_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_113_nl = MUX_v_64_2_2(input_mem_banks_bank_a_56_sva_dfm_2,
      input_mem_banks_bank_a_56_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_115_nl = MUX_v_64_2_2(input_mem_banks_bank_a_57_sva_dfm_2,
      input_mem_banks_bank_a_57_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_117_nl = MUX_v_64_2_2(input_mem_banks_bank_a_58_sva_dfm_2,
      input_mem_banks_bank_a_58_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_119_nl = MUX_v_64_2_2(input_mem_banks_bank_a_59_sva_dfm_2,
      input_mem_banks_bank_a_59_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_121_nl = MUX_v_64_2_2(input_mem_banks_bank_a_60_sva_dfm_2,
      input_mem_banks_bank_a_60_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_123_nl = MUX_v_64_2_2(input_mem_banks_bank_a_61_sva_dfm_2,
      input_mem_banks_bank_a_61_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_125_nl = MUX_v_64_2_2(input_mem_banks_bank_a_62_sva_dfm_2,
      input_mem_banks_bank_a_62_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_127_nl = MUX_v_64_2_2(input_mem_banks_bank_a_63_sva_dfm_2,
      input_mem_banks_bank_a_63_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_129_nl = MUX_v_64_2_2(input_mem_banks_bank_a_64_sva_dfm_2,
      input_mem_banks_bank_a_64_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_131_nl = MUX_v_64_2_2(input_mem_banks_bank_a_65_sva_dfm_2,
      input_mem_banks_bank_a_65_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_133_nl = MUX_v_64_2_2(input_mem_banks_bank_a_66_sva_dfm_2,
      input_mem_banks_bank_a_66_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_135_nl = MUX_v_64_2_2(input_mem_banks_bank_a_67_sva_dfm_2,
      input_mem_banks_bank_a_67_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_137_nl = MUX_v_64_2_2(input_mem_banks_bank_a_68_sva_dfm_2,
      input_mem_banks_bank_a_68_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_139_nl = MUX_v_64_2_2(input_mem_banks_bank_a_69_sva_dfm_2,
      input_mem_banks_bank_a_69_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_141_nl = MUX_v_64_2_2(input_mem_banks_bank_a_70_sva_dfm_2,
      input_mem_banks_bank_a_70_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_143_nl = MUX_v_64_2_2(input_mem_banks_bank_a_71_sva_dfm_2,
      input_mem_banks_bank_a_71_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_145_nl = MUX_v_64_2_2(input_mem_banks_bank_a_72_sva_dfm_2,
      input_mem_banks_bank_a_72_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_147_nl = MUX_v_64_2_2(input_mem_banks_bank_a_73_sva_dfm_2,
      input_mem_banks_bank_a_73_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_149_nl = MUX_v_64_2_2(input_mem_banks_bank_a_74_sva_dfm_2,
      input_mem_banks_bank_a_74_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_151_nl = MUX_v_64_2_2(input_mem_banks_bank_a_75_sva_dfm_2,
      input_mem_banks_bank_a_75_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_153_nl = MUX_v_64_2_2(input_mem_banks_bank_a_76_sva_dfm_2,
      input_mem_banks_bank_a_76_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_155_nl = MUX_v_64_2_2(input_mem_banks_bank_a_77_sva_dfm_2,
      input_mem_banks_bank_a_77_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_157_nl = MUX_v_64_2_2(input_mem_banks_bank_a_78_sva_dfm_2,
      input_mem_banks_bank_a_78_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_159_nl = MUX_v_64_2_2(input_mem_banks_bank_a_79_sva_dfm_2,
      input_mem_banks_bank_a_79_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_161_nl = MUX_v_64_2_2(input_mem_banks_bank_a_80_sva_dfm_2,
      input_mem_banks_bank_a_80_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_163_nl = MUX_v_64_2_2(input_mem_banks_bank_a_81_sva_dfm_2,
      input_mem_banks_bank_a_81_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_165_nl = MUX_v_64_2_2(input_mem_banks_bank_a_82_sva_dfm_2,
      input_mem_banks_bank_a_82_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_167_nl = MUX_v_64_2_2(input_mem_banks_bank_a_83_sva_dfm_2,
      input_mem_banks_bank_a_83_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_169_nl = MUX_v_64_2_2(input_mem_banks_bank_a_84_sva_dfm_2,
      input_mem_banks_bank_a_84_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_171_nl = MUX_v_64_2_2(input_mem_banks_bank_a_85_sva_dfm_2,
      input_mem_banks_bank_a_85_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_173_nl = MUX_v_64_2_2(input_mem_banks_bank_a_86_sva_dfm_2,
      input_mem_banks_bank_a_86_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_175_nl = MUX_v_64_2_2(input_mem_banks_bank_a_87_sva_dfm_2,
      input_mem_banks_bank_a_87_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_177_nl = MUX_v_64_2_2(input_mem_banks_bank_a_88_sva_dfm_2,
      input_mem_banks_bank_a_88_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_179_nl = MUX_v_64_2_2(input_mem_banks_bank_a_89_sva_dfm_2,
      input_mem_banks_bank_a_89_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_181_nl = MUX_v_64_2_2(input_mem_banks_bank_a_90_sva_dfm_2,
      input_mem_banks_bank_a_90_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_183_nl = MUX_v_64_2_2(input_mem_banks_bank_a_91_sva_dfm_2,
      input_mem_banks_bank_a_91_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_185_nl = MUX_v_64_2_2(input_mem_banks_bank_a_92_sva_dfm_2,
      input_mem_banks_bank_a_92_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_187_nl = MUX_v_64_2_2(input_mem_banks_bank_a_93_sva_dfm_2,
      input_mem_banks_bank_a_93_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_189_nl = MUX_v_64_2_2(input_mem_banks_bank_a_94_sva_dfm_2,
      input_mem_banks_bank_a_94_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_191_nl = MUX_v_64_2_2(input_mem_banks_bank_a_95_sva_dfm_2,
      input_mem_banks_bank_a_95_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_193_nl = MUX_v_64_2_2(input_mem_banks_bank_a_96_sva_dfm_2,
      input_mem_banks_bank_a_96_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_195_nl = MUX_v_64_2_2(input_mem_banks_bank_a_97_sva_dfm_2,
      input_mem_banks_bank_a_97_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_197_nl = MUX_v_64_2_2(input_mem_banks_bank_a_98_sva_dfm_2,
      input_mem_banks_bank_a_98_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_199_nl = MUX_v_64_2_2(input_mem_banks_bank_a_99_sva_dfm_2,
      input_mem_banks_bank_a_99_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_201_nl = MUX_v_64_2_2(input_mem_banks_bank_a_100_sva_dfm_2,
      input_mem_banks_bank_a_100_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_203_nl = MUX_v_64_2_2(input_mem_banks_bank_a_101_sva_dfm_2,
      input_mem_banks_bank_a_101_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_205_nl = MUX_v_64_2_2(input_mem_banks_bank_a_102_sva_dfm_2,
      input_mem_banks_bank_a_102_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_207_nl = MUX_v_64_2_2(input_mem_banks_bank_a_103_sva_dfm_2,
      input_mem_banks_bank_a_103_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_209_nl = MUX_v_64_2_2(input_mem_banks_bank_a_104_sva_dfm_2,
      input_mem_banks_bank_a_104_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_211_nl = MUX_v_64_2_2(input_mem_banks_bank_a_105_sva_dfm_2,
      input_mem_banks_bank_a_105_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_213_nl = MUX_v_64_2_2(input_mem_banks_bank_a_106_sva_dfm_2,
      input_mem_banks_bank_a_106_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_215_nl = MUX_v_64_2_2(input_mem_banks_bank_a_107_sva_dfm_2,
      input_mem_banks_bank_a_107_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_217_nl = MUX_v_64_2_2(input_mem_banks_bank_a_108_sva_dfm_2,
      input_mem_banks_bank_a_108_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_219_nl = MUX_v_64_2_2(input_mem_banks_bank_a_109_sva_dfm_2,
      input_mem_banks_bank_a_109_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_221_nl = MUX_v_64_2_2(input_mem_banks_bank_a_110_sva_dfm_2,
      input_mem_banks_bank_a_110_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_223_nl = MUX_v_64_2_2(input_mem_banks_bank_a_111_sva_dfm_2,
      input_mem_banks_bank_a_111_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_225_nl = MUX_v_64_2_2(input_mem_banks_bank_a_112_sva_dfm_2,
      input_mem_banks_bank_a_112_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_227_nl = MUX_v_64_2_2(input_mem_banks_bank_a_113_sva_dfm_2,
      input_mem_banks_bank_a_113_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_229_nl = MUX_v_64_2_2(input_mem_banks_bank_a_114_sva_dfm_2,
      input_mem_banks_bank_a_114_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_231_nl = MUX_v_64_2_2(input_mem_banks_bank_a_115_sva_dfm_2,
      input_mem_banks_bank_a_115_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_233_nl = MUX_v_64_2_2(input_mem_banks_bank_a_116_sva_dfm_2,
      input_mem_banks_bank_a_116_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_235_nl = MUX_v_64_2_2(input_mem_banks_bank_a_117_sva_dfm_2,
      input_mem_banks_bank_a_117_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_237_nl = MUX_v_64_2_2(input_mem_banks_bank_a_118_sva_dfm_2,
      input_mem_banks_bank_a_118_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_239_nl = MUX_v_64_2_2(input_mem_banks_bank_a_119_sva_dfm_2,
      input_mem_banks_bank_a_119_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_241_nl = MUX_v_64_2_2(input_mem_banks_bank_a_120_sva_dfm_2,
      input_mem_banks_bank_a_120_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_243_nl = MUX_v_64_2_2(input_mem_banks_bank_a_121_sva_dfm_2,
      input_mem_banks_bank_a_121_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_245_nl = MUX_v_64_2_2(input_mem_banks_bank_a_122_sva_dfm_2,
      input_mem_banks_bank_a_122_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_247_nl = MUX_v_64_2_2(input_mem_banks_bank_a_123_sva_dfm_2,
      input_mem_banks_bank_a_123_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_249_nl = MUX_v_64_2_2(input_mem_banks_bank_a_124_sva_dfm_2,
      input_mem_banks_bank_a_124_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_251_nl = MUX_v_64_2_2(input_mem_banks_bank_a_125_sva_dfm_2,
      input_mem_banks_bank_a_125_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_253_nl = MUX_v_64_2_2(input_mem_banks_bank_a_126_sva_dfm_2,
      input_mem_banks_bank_a_126_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_255_nl = MUX_v_64_2_2(input_mem_banks_bank_a_127_sva_dfm_2,
      input_mem_banks_bank_a_127_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_257_nl = MUX_v_64_2_2(input_mem_banks_bank_a_128_sva_dfm_2,
      input_mem_banks_bank_a_128_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_259_nl = MUX_v_64_2_2(input_mem_banks_bank_a_129_sva_dfm_2,
      input_mem_banks_bank_a_129_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_261_nl = MUX_v_64_2_2(input_mem_banks_bank_a_130_sva_dfm_2,
      input_mem_banks_bank_a_130_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_263_nl = MUX_v_64_2_2(input_mem_banks_bank_a_131_sva_dfm_2,
      input_mem_banks_bank_a_131_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_265_nl = MUX_v_64_2_2(input_mem_banks_bank_a_132_sva_dfm_2,
      input_mem_banks_bank_a_132_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_267_nl = MUX_v_64_2_2(input_mem_banks_bank_a_133_sva_dfm_2,
      input_mem_banks_bank_a_133_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_269_nl = MUX_v_64_2_2(input_mem_banks_bank_a_134_sva_dfm_2,
      input_mem_banks_bank_a_134_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_271_nl = MUX_v_64_2_2(input_mem_banks_bank_a_135_sva_dfm_2,
      input_mem_banks_bank_a_135_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_273_nl = MUX_v_64_2_2(input_mem_banks_bank_a_136_sva_dfm_2,
      input_mem_banks_bank_a_136_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_275_nl = MUX_v_64_2_2(input_mem_banks_bank_a_137_sva_dfm_2,
      input_mem_banks_bank_a_137_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_277_nl = MUX_v_64_2_2(input_mem_banks_bank_a_138_sva_dfm_2,
      input_mem_banks_bank_a_138_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_279_nl = MUX_v_64_2_2(input_mem_banks_bank_a_139_sva_dfm_2,
      input_mem_banks_bank_a_139_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_281_nl = MUX_v_64_2_2(input_mem_banks_bank_a_140_sva_dfm_2,
      input_mem_banks_bank_a_140_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_283_nl = MUX_v_64_2_2(input_mem_banks_bank_a_141_sva_dfm_2,
      input_mem_banks_bank_a_141_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_285_nl = MUX_v_64_2_2(input_mem_banks_bank_a_142_sva_dfm_2,
      input_mem_banks_bank_a_142_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_287_nl = MUX_v_64_2_2(input_mem_banks_bank_a_143_sva_dfm_2,
      input_mem_banks_bank_a_143_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_289_nl = MUX_v_64_2_2(input_mem_banks_bank_a_144_sva_dfm_2,
      input_mem_banks_bank_a_144_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_291_nl = MUX_v_64_2_2(input_mem_banks_bank_a_145_sva_dfm_2,
      input_mem_banks_bank_a_145_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_293_nl = MUX_v_64_2_2(input_mem_banks_bank_a_146_sva_dfm_2,
      input_mem_banks_bank_a_146_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_295_nl = MUX_v_64_2_2(input_mem_banks_bank_a_147_sva_dfm_2,
      input_mem_banks_bank_a_147_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_297_nl = MUX_v_64_2_2(input_mem_banks_bank_a_148_sva_dfm_2,
      input_mem_banks_bank_a_148_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_299_nl = MUX_v_64_2_2(input_mem_banks_bank_a_149_sva_dfm_2,
      input_mem_banks_bank_a_149_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_301_nl = MUX_v_64_2_2(input_mem_banks_bank_a_150_sva_dfm_2,
      input_mem_banks_bank_a_150_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_303_nl = MUX_v_64_2_2(input_mem_banks_bank_a_151_sva_dfm_2,
      input_mem_banks_bank_a_151_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_305_nl = MUX_v_64_2_2(input_mem_banks_bank_a_152_sva_dfm_2,
      input_mem_banks_bank_a_152_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_307_nl = MUX_v_64_2_2(input_mem_banks_bank_a_153_sva_dfm_2,
      input_mem_banks_bank_a_153_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_309_nl = MUX_v_64_2_2(input_mem_banks_bank_a_154_sva_dfm_2,
      input_mem_banks_bank_a_154_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_311_nl = MUX_v_64_2_2(input_mem_banks_bank_a_155_sva_dfm_2,
      input_mem_banks_bank_a_155_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_313_nl = MUX_v_64_2_2(input_mem_banks_bank_a_156_sva_dfm_2,
      input_mem_banks_bank_a_156_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_315_nl = MUX_v_64_2_2(input_mem_banks_bank_a_157_sva_dfm_2,
      input_mem_banks_bank_a_157_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_317_nl = MUX_v_64_2_2(input_mem_banks_bank_a_158_sva_dfm_2,
      input_mem_banks_bank_a_158_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_319_nl = MUX_v_64_2_2(input_mem_banks_bank_a_159_sva_dfm_2,
      input_mem_banks_bank_a_159_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_321_nl = MUX_v_64_2_2(input_mem_banks_bank_a_160_sva_dfm_2,
      input_mem_banks_bank_a_160_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_323_nl = MUX_v_64_2_2(input_mem_banks_bank_a_161_sva_dfm_2,
      input_mem_banks_bank_a_161_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_325_nl = MUX_v_64_2_2(input_mem_banks_bank_a_162_sva_dfm_2,
      input_mem_banks_bank_a_162_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_327_nl = MUX_v_64_2_2(input_mem_banks_bank_a_163_sva_dfm_2,
      input_mem_banks_bank_a_163_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_329_nl = MUX_v_64_2_2(input_mem_banks_bank_a_164_sva_dfm_2,
      input_mem_banks_bank_a_164_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_331_nl = MUX_v_64_2_2(input_mem_banks_bank_a_165_sva_dfm_2,
      input_mem_banks_bank_a_165_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_333_nl = MUX_v_64_2_2(input_mem_banks_bank_a_166_sva_dfm_2,
      input_mem_banks_bank_a_166_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_335_nl = MUX_v_64_2_2(input_mem_banks_bank_a_167_sva_dfm_2,
      input_mem_banks_bank_a_167_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_337_nl = MUX_v_64_2_2(input_mem_banks_bank_a_168_sva_dfm_2,
      input_mem_banks_bank_a_168_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_339_nl = MUX_v_64_2_2(input_mem_banks_bank_a_169_sva_dfm_2,
      input_mem_banks_bank_a_169_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_341_nl = MUX_v_64_2_2(input_mem_banks_bank_a_170_sva_dfm_2,
      input_mem_banks_bank_a_170_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_343_nl = MUX_v_64_2_2(input_mem_banks_bank_a_171_sva_dfm_2,
      input_mem_banks_bank_a_171_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_345_nl = MUX_v_64_2_2(input_mem_banks_bank_a_172_sva_dfm_2,
      input_mem_banks_bank_a_172_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_347_nl = MUX_v_64_2_2(input_mem_banks_bank_a_173_sva_dfm_2,
      input_mem_banks_bank_a_173_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_349_nl = MUX_v_64_2_2(input_mem_banks_bank_a_174_sva_dfm_2,
      input_mem_banks_bank_a_174_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_351_nl = MUX_v_64_2_2(input_mem_banks_bank_a_175_sva_dfm_2,
      input_mem_banks_bank_a_175_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_353_nl = MUX_v_64_2_2(input_mem_banks_bank_a_176_sva_dfm_2,
      input_mem_banks_bank_a_176_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_355_nl = MUX_v_64_2_2(input_mem_banks_bank_a_177_sva_dfm_2,
      input_mem_banks_bank_a_177_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_357_nl = MUX_v_64_2_2(input_mem_banks_bank_a_178_sva_dfm_2,
      input_mem_banks_bank_a_178_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_359_nl = MUX_v_64_2_2(input_mem_banks_bank_a_179_sva_dfm_2,
      input_mem_banks_bank_a_179_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_361_nl = MUX_v_64_2_2(input_mem_banks_bank_a_180_sva_dfm_2,
      input_mem_banks_bank_a_180_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_363_nl = MUX_v_64_2_2(input_mem_banks_bank_a_181_sva_dfm_2,
      input_mem_banks_bank_a_181_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_365_nl = MUX_v_64_2_2(input_mem_banks_bank_a_182_sva_dfm_2,
      input_mem_banks_bank_a_182_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_367_nl = MUX_v_64_2_2(input_mem_banks_bank_a_183_sva_dfm_2,
      input_mem_banks_bank_a_183_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_369_nl = MUX_v_64_2_2(input_mem_banks_bank_a_184_sva_dfm_2,
      input_mem_banks_bank_a_184_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_371_nl = MUX_v_64_2_2(input_mem_banks_bank_a_185_sva_dfm_2,
      input_mem_banks_bank_a_185_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_373_nl = MUX_v_64_2_2(input_mem_banks_bank_a_186_sva_dfm_2,
      input_mem_banks_bank_a_186_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_375_nl = MUX_v_64_2_2(input_mem_banks_bank_a_187_sva_dfm_2,
      input_mem_banks_bank_a_187_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_377_nl = MUX_v_64_2_2(input_mem_banks_bank_a_188_sva_dfm_2,
      input_mem_banks_bank_a_188_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_379_nl = MUX_v_64_2_2(input_mem_banks_bank_a_189_sva_dfm_2,
      input_mem_banks_bank_a_189_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_381_nl = MUX_v_64_2_2(input_mem_banks_bank_a_190_sva_dfm_2,
      input_mem_banks_bank_a_190_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_383_nl = MUX_v_64_2_2(input_mem_banks_bank_a_191_sva_dfm_2,
      input_mem_banks_bank_a_191_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_385_nl = MUX_v_64_2_2(input_mem_banks_bank_a_192_sva_dfm_2,
      input_mem_banks_bank_a_192_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_387_nl = MUX_v_64_2_2(input_mem_banks_bank_a_193_sva_dfm_2,
      input_mem_banks_bank_a_193_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_389_nl = MUX_v_64_2_2(input_mem_banks_bank_a_194_sva_dfm_2,
      input_mem_banks_bank_a_194_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_391_nl = MUX_v_64_2_2(input_mem_banks_bank_a_195_sva_dfm_2,
      input_mem_banks_bank_a_195_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_393_nl = MUX_v_64_2_2(input_mem_banks_bank_a_196_sva_dfm_2,
      input_mem_banks_bank_a_196_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_395_nl = MUX_v_64_2_2(input_mem_banks_bank_a_197_sva_dfm_2,
      input_mem_banks_bank_a_197_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_397_nl = MUX_v_64_2_2(input_mem_banks_bank_a_198_sva_dfm_2,
      input_mem_banks_bank_a_198_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_399_nl = MUX_v_64_2_2(input_mem_banks_bank_a_199_sva_dfm_2,
      input_mem_banks_bank_a_199_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_401_nl = MUX_v_64_2_2(input_mem_banks_bank_a_200_sva_dfm_2,
      input_mem_banks_bank_a_200_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_403_nl = MUX_v_64_2_2(input_mem_banks_bank_a_201_sva_dfm_2,
      input_mem_banks_bank_a_201_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_405_nl = MUX_v_64_2_2(input_mem_banks_bank_a_202_sva_dfm_2,
      input_mem_banks_bank_a_202_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_407_nl = MUX_v_64_2_2(input_mem_banks_bank_a_203_sva_dfm_2,
      input_mem_banks_bank_a_203_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_409_nl = MUX_v_64_2_2(input_mem_banks_bank_a_204_sva_dfm_2,
      input_mem_banks_bank_a_204_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_411_nl = MUX_v_64_2_2(input_mem_banks_bank_a_205_sva_dfm_2,
      input_mem_banks_bank_a_205_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_413_nl = MUX_v_64_2_2(input_mem_banks_bank_a_206_sva_dfm_2,
      input_mem_banks_bank_a_206_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_415_nl = MUX_v_64_2_2(input_mem_banks_bank_a_207_sva_dfm_2,
      input_mem_banks_bank_a_207_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_417_nl = MUX_v_64_2_2(input_mem_banks_bank_a_208_sva_dfm_2,
      input_mem_banks_bank_a_208_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_419_nl = MUX_v_64_2_2(input_mem_banks_bank_a_209_sva_dfm_2,
      input_mem_banks_bank_a_209_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_421_nl = MUX_v_64_2_2(input_mem_banks_bank_a_210_sva_dfm_2,
      input_mem_banks_bank_a_210_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_423_nl = MUX_v_64_2_2(input_mem_banks_bank_a_211_sva_dfm_2,
      input_mem_banks_bank_a_211_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_425_nl = MUX_v_64_2_2(input_mem_banks_bank_a_212_sva_dfm_2,
      input_mem_banks_bank_a_212_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_427_nl = MUX_v_64_2_2(input_mem_banks_bank_a_213_sva_dfm_2,
      input_mem_banks_bank_a_213_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_429_nl = MUX_v_64_2_2(input_mem_banks_bank_a_214_sva_dfm_2,
      input_mem_banks_bank_a_214_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_431_nl = MUX_v_64_2_2(input_mem_banks_bank_a_215_sva_dfm_2,
      input_mem_banks_bank_a_215_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_433_nl = MUX_v_64_2_2(input_mem_banks_bank_a_216_sva_dfm_2,
      input_mem_banks_bank_a_216_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_435_nl = MUX_v_64_2_2(input_mem_banks_bank_a_217_sva_dfm_2,
      input_mem_banks_bank_a_217_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_437_nl = MUX_v_64_2_2(input_mem_banks_bank_a_218_sva_dfm_2,
      input_mem_banks_bank_a_218_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_439_nl = MUX_v_64_2_2(input_mem_banks_bank_a_219_sva_dfm_2,
      input_mem_banks_bank_a_219_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_441_nl = MUX_v_64_2_2(input_mem_banks_bank_a_220_sva_dfm_2,
      input_mem_banks_bank_a_220_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_443_nl = MUX_v_64_2_2(input_mem_banks_bank_a_221_sva_dfm_2,
      input_mem_banks_bank_a_221_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_445_nl = MUX_v_64_2_2(input_mem_banks_bank_a_222_sva_dfm_2,
      input_mem_banks_bank_a_222_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_447_nl = MUX_v_64_2_2(input_mem_banks_bank_a_223_sva_dfm_2,
      input_mem_banks_bank_a_223_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_449_nl = MUX_v_64_2_2(input_mem_banks_bank_a_224_sva_dfm_2,
      input_mem_banks_bank_a_224_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_451_nl = MUX_v_64_2_2(input_mem_banks_bank_a_225_sva_dfm_2,
      input_mem_banks_bank_a_225_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_453_nl = MUX_v_64_2_2(input_mem_banks_bank_a_226_sva_dfm_2,
      input_mem_banks_bank_a_226_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_455_nl = MUX_v_64_2_2(input_mem_banks_bank_a_227_sva_dfm_2,
      input_mem_banks_bank_a_227_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_457_nl = MUX_v_64_2_2(input_mem_banks_bank_a_228_sva_dfm_2,
      input_mem_banks_bank_a_228_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_459_nl = MUX_v_64_2_2(input_mem_banks_bank_a_229_sva_dfm_2,
      input_mem_banks_bank_a_229_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_461_nl = MUX_v_64_2_2(input_mem_banks_bank_a_230_sva_dfm_2,
      input_mem_banks_bank_a_230_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_463_nl = MUX_v_64_2_2(input_mem_banks_bank_a_231_sva_dfm_2,
      input_mem_banks_bank_a_231_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_465_nl = MUX_v_64_2_2(input_mem_banks_bank_a_232_sva_dfm_2,
      input_mem_banks_bank_a_232_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_467_nl = MUX_v_64_2_2(input_mem_banks_bank_a_233_sva_dfm_2,
      input_mem_banks_bank_a_233_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_469_nl = MUX_v_64_2_2(input_mem_banks_bank_a_234_sva_dfm_2,
      input_mem_banks_bank_a_234_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_471_nl = MUX_v_64_2_2(input_mem_banks_bank_a_235_sva_dfm_2,
      input_mem_banks_bank_a_235_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_473_nl = MUX_v_64_2_2(input_mem_banks_bank_a_236_sva_dfm_2,
      input_mem_banks_bank_a_236_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_475_nl = MUX_v_64_2_2(input_mem_banks_bank_a_237_sva_dfm_2,
      input_mem_banks_bank_a_237_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_477_nl = MUX_v_64_2_2(input_mem_banks_bank_a_238_sva_dfm_2,
      input_mem_banks_bank_a_238_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_479_nl = MUX_v_64_2_2(input_mem_banks_bank_a_239_sva_dfm_2,
      input_mem_banks_bank_a_239_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_481_nl = MUX_v_64_2_2(input_mem_banks_bank_a_240_sva_dfm_2,
      input_mem_banks_bank_a_240_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_483_nl = MUX_v_64_2_2(input_mem_banks_bank_a_241_sva_dfm_2,
      input_mem_banks_bank_a_241_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_485_nl = MUX_v_64_2_2(input_mem_banks_bank_a_242_sva_dfm_2,
      input_mem_banks_bank_a_242_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_487_nl = MUX_v_64_2_2(input_mem_banks_bank_a_243_sva_dfm_2,
      input_mem_banks_bank_a_243_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_489_nl = MUX_v_64_2_2(input_mem_banks_bank_a_244_sva_dfm_2,
      input_mem_banks_bank_a_244_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_491_nl = MUX_v_64_2_2(input_mem_banks_bank_a_245_sva_dfm_2,
      input_mem_banks_bank_a_245_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_493_nl = MUX_v_64_2_2(input_mem_banks_bank_a_246_sva_dfm_2,
      input_mem_banks_bank_a_246_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_495_nl = MUX_v_64_2_2(input_mem_banks_bank_a_247_sva_dfm_2,
      input_mem_banks_bank_a_247_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_497_nl = MUX_v_64_2_2(input_mem_banks_bank_a_248_sva_dfm_2,
      input_mem_banks_bank_a_248_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_499_nl = MUX_v_64_2_2(input_mem_banks_bank_a_249_sva_dfm_2,
      input_mem_banks_bank_a_249_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_501_nl = MUX_v_64_2_2(input_mem_banks_bank_a_250_sva_dfm_2,
      input_mem_banks_bank_a_250_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_503_nl = MUX_v_64_2_2(input_mem_banks_bank_a_251_sva_dfm_2,
      input_mem_banks_bank_a_251_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_505_nl = MUX_v_64_2_2(input_mem_banks_bank_a_252_sva_dfm_2,
      input_mem_banks_bank_a_252_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_507_nl = MUX_v_64_2_2(input_mem_banks_bank_a_253_sva_dfm_2,
      input_mem_banks_bank_a_253_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_509_nl = MUX_v_64_2_2(input_mem_banks_bank_a_254_sva_dfm_2,
      input_mem_banks_bank_a_254_sva_dfm_2_mx0w0, while_stage_0_3);
  assign input_mem_banks_bank_a_mux_511_nl = MUX_v_64_2_2(input_mem_banks_bank_a_255_sva_dfm_2,
      input_mem_banks_bank_a_255_sva_dfm_2_mx0w0, while_stage_0_3);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl = MUX_v_4_2_2(pe_config_num_manager_sva,
      (pe_manager_base_bias_sva[3:0]), and_301_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl = MUX_v_7_2_2((pe_config_num_output_sva[6:0]),
      (pe_manager_base_bias_sva[14:8]), and_301_cse);
  assign weight_mem_banks_load_store_for_else_mux1h_8_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[63]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[39]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[39]),
      {and_dcpl_594 , and_dcpl_595 , and_dcpl_597});
  assign weight_mem_banks_load_store_for_else_mux1h_38_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[62:56]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[38:32]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[38:32]),
      rva_out_reg_data_46_40_sva_dfm_1_4, {and_dcpl_594 , and_dcpl_595 , and_dcpl_597
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2208_nl = ~ or_dcpl_297;
  assign weight_mem_banks_load_store_for_else_mux1h_15_nl = MUX1HOT_v_4_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[47:44]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[31:28]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[31:28]),
      {and_dcpl_594 , and_dcpl_595 , and_dcpl_597});
  assign not_2209_nl = ~ or_dcpl_297;
  assign weight_mem_banks_load_store_for_else_mux1h_39_nl = MUX1HOT_v_4_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[43:40]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[27:24]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[27:24]),
      rva_out_reg_data_35_32_sva_dfm_1_4, {and_dcpl_594 , and_dcpl_595 , and_dcpl_597
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2210_nl = ~ or_dcpl_297;
  assign weight_mem_banks_load_store_for_else_mux1h_22_nl = MUX1HOT_v_2_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[39:38]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[23:22]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[23:22]),
      {and_dcpl_594 , and_dcpl_595 , and_dcpl_597});
  assign not_2211_nl = ~ or_dcpl_297;
  assign weight_mem_banks_load_store_for_else_mux1h_40_nl = MUX1HOT_v_6_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[37:32]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[21:16]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[21:16]),
      rva_out_reg_data_30_25_sva_dfm_2, {and_dcpl_594 , and_dcpl_595 , and_dcpl_597
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2212_nl = ~ or_dcpl_297;
  assign weight_mem_banks_load_store_for_else_mux1h_27_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[31]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[15]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[15]),
      {and_dcpl_594 , and_dcpl_595 , and_dcpl_597});
  assign weight_mem_banks_load_store_for_else_mux1h_41_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[30:24]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[14:8]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[14:8]),
      rva_out_reg_data_23_17_sva_dfm_2, {and_dcpl_594 , and_dcpl_595 , and_dcpl_597
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2214_nl = ~ or_dcpl_297;
  assign weight_mem_banks_load_store_for_else_mux1h_32_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[23]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[7]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[7]),
      {and_dcpl_594 , and_dcpl_595 , and_dcpl_597});
  assign weight_mem_banks_load_store_for_else_mux1h_42_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[22:16]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[6:0]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[6:0]),
      rva_out_reg_data_15_9_sva_dfm_4, {and_dcpl_594 , and_dcpl_595 , and_dcpl_597
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2216_nl = ~ or_dcpl_297;
  assign and_2185_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2
      | reg_weight_mem_run_3_for_5_and_165_itm_2_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2
      | reg_weight_mem_run_3_for_5_and_163_itm_2_cse | reg_weight_mem_run_3_for_5_and_162_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign mux_887_nl = MUX_s_1_2_2(and_2185_nl, or_2320_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_2188_nl = (reg_weight_mem_run_3_for_5_and_168_itm_2_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2 | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_162_itm_2_cse | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign or_2341_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1 | and_1840_cse;
  assign mux_896_nl = MUX_s_1_2_2(and_2188_nl, or_2341_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_2189_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2
      | reg_weight_mem_run_3_for_5_and_167_itm_2_cse | reg_weight_mem_run_3_for_5_and_166_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_165_itm_2_cse | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2
      | reg_weight_mem_run_3_for_5_and_163_itm_2_cse | reg_weight_mem_run_3_for_5_and_162_itm_2_cse
      | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse) & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign mux_899_nl = MUX_s_1_2_2(and_2189_nl, or_2320_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_2355_nl = or_tmp_1863 | and_1831_cse;
  assign mux_902_nl = MUX_s_1_2_2(and_2190_cse, or_2355_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_905_nl = MUX_s_1_2_2(and_2190_cse, or_2320_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_2371_nl = reg_weight_mem_run_3_for_5_and_168_itm_2_cse | reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_166_itm_2_cse | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | weight_mem_run_3_for_5_and_164_itm_2 | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_162_itm_2_cse | weight_mem_run_3_for_5_and_182_cse;
  assign or_2369_nl = or_tmp_1863 | and_1840_cse;
  assign mux_908_nl = MUX_s_1_2_2(or_2371_nl, or_2369_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_9_2;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [8:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_8_2;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [7:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    result = result | (input_5 & {11{sel[5]}});
    result = result | (input_6 & {11{sel[6]}});
    result = result | (input_7 & {11{sel[7]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_8_2;
    input [2:0] input_7;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [7:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    result = result | (input_6 & {3{sel[6]}});
    result = result | (input_7 & {3{sel[7]}});
    MUX1HOT_v_3_8_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_9_2;
    input [2:0] input_8;
    input [2:0] input_7;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [8:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    result = result | (input_6 & {3{sel[6]}});
    result = result | (input_7 & {3{sel[7]}});
    result = result | (input_8 & {3{sel[8]}});
    MUX1HOT_v_3_9_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_8_2;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [7:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    MUX1HOT_v_4_8_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_9_2;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [8:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    MUX1HOT_v_4_9_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | (input_1 & {64{sel[1]}});
    result = result | (input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_8_2;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [7:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    MUX1HOT_v_6_8_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_9_2;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [8:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    result = result | (input_8 & {6{sel[8]}});
    MUX1HOT_v_6_9_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_8_2;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [7:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    result = result | (input_6 & {7{sel[6]}});
    result = result | (input_7 & {7{sel[7]}});
    MUX1HOT_v_7_8_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_9_2;
    input [6:0] input_8;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [8:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    result = result | (input_6 & {7{sel[6]}});
    result = result | (input_7 & {7{sel[7]}});
    result = result | (input_8 & {7{sel[8]}});
    MUX1HOT_v_7_9_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_5_2;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [4:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    MUX1HOT_v_8_5_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_8_2;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [7:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    MUX1HOT_v_8_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_9_2;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [8:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    result = result | (input_8 & {8{sel[8]}});
    MUX1HOT_v_8_9_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_8_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input [2:0] sel;
    reg  result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_s_1_8_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_8_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [10:0] input_2;
    input [10:0] input_3;
    input [10:0] input_4;
    input [10:0] input_5;
    input [10:0] input_6;
    input [10:0] input_7;
    input [2:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_11_8_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input  sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input  sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [18:0] MUX_v_19_2_2;
    input [18:0] input_0;
    input [18:0] input_1;
    input  sel;
    reg [18:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_19_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_8_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [2:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_4_8_2 = result;
  end
  endfunction


  function automatic [55:0] MUX_v_56_2_2;
    input [55:0] input_0;
    input [55:0] input_1;
    input  sel;
    reg [55:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_56_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_256_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [63:0] input_2;
    input [63:0] input_3;
    input [63:0] input_4;
    input [63:0] input_5;
    input [63:0] input_6;
    input [63:0] input_7;
    input [63:0] input_8;
    input [63:0] input_9;
    input [63:0] input_10;
    input [63:0] input_11;
    input [63:0] input_12;
    input [63:0] input_13;
    input [63:0] input_14;
    input [63:0] input_15;
    input [63:0] input_16;
    input [63:0] input_17;
    input [63:0] input_18;
    input [63:0] input_19;
    input [63:0] input_20;
    input [63:0] input_21;
    input [63:0] input_22;
    input [63:0] input_23;
    input [63:0] input_24;
    input [63:0] input_25;
    input [63:0] input_26;
    input [63:0] input_27;
    input [63:0] input_28;
    input [63:0] input_29;
    input [63:0] input_30;
    input [63:0] input_31;
    input [63:0] input_32;
    input [63:0] input_33;
    input [63:0] input_34;
    input [63:0] input_35;
    input [63:0] input_36;
    input [63:0] input_37;
    input [63:0] input_38;
    input [63:0] input_39;
    input [63:0] input_40;
    input [63:0] input_41;
    input [63:0] input_42;
    input [63:0] input_43;
    input [63:0] input_44;
    input [63:0] input_45;
    input [63:0] input_46;
    input [63:0] input_47;
    input [63:0] input_48;
    input [63:0] input_49;
    input [63:0] input_50;
    input [63:0] input_51;
    input [63:0] input_52;
    input [63:0] input_53;
    input [63:0] input_54;
    input [63:0] input_55;
    input [63:0] input_56;
    input [63:0] input_57;
    input [63:0] input_58;
    input [63:0] input_59;
    input [63:0] input_60;
    input [63:0] input_61;
    input [63:0] input_62;
    input [63:0] input_63;
    input [63:0] input_64;
    input [63:0] input_65;
    input [63:0] input_66;
    input [63:0] input_67;
    input [63:0] input_68;
    input [63:0] input_69;
    input [63:0] input_70;
    input [63:0] input_71;
    input [63:0] input_72;
    input [63:0] input_73;
    input [63:0] input_74;
    input [63:0] input_75;
    input [63:0] input_76;
    input [63:0] input_77;
    input [63:0] input_78;
    input [63:0] input_79;
    input [63:0] input_80;
    input [63:0] input_81;
    input [63:0] input_82;
    input [63:0] input_83;
    input [63:0] input_84;
    input [63:0] input_85;
    input [63:0] input_86;
    input [63:0] input_87;
    input [63:0] input_88;
    input [63:0] input_89;
    input [63:0] input_90;
    input [63:0] input_91;
    input [63:0] input_92;
    input [63:0] input_93;
    input [63:0] input_94;
    input [63:0] input_95;
    input [63:0] input_96;
    input [63:0] input_97;
    input [63:0] input_98;
    input [63:0] input_99;
    input [63:0] input_100;
    input [63:0] input_101;
    input [63:0] input_102;
    input [63:0] input_103;
    input [63:0] input_104;
    input [63:0] input_105;
    input [63:0] input_106;
    input [63:0] input_107;
    input [63:0] input_108;
    input [63:0] input_109;
    input [63:0] input_110;
    input [63:0] input_111;
    input [63:0] input_112;
    input [63:0] input_113;
    input [63:0] input_114;
    input [63:0] input_115;
    input [63:0] input_116;
    input [63:0] input_117;
    input [63:0] input_118;
    input [63:0] input_119;
    input [63:0] input_120;
    input [63:0] input_121;
    input [63:0] input_122;
    input [63:0] input_123;
    input [63:0] input_124;
    input [63:0] input_125;
    input [63:0] input_126;
    input [63:0] input_127;
    input [63:0] input_128;
    input [63:0] input_129;
    input [63:0] input_130;
    input [63:0] input_131;
    input [63:0] input_132;
    input [63:0] input_133;
    input [63:0] input_134;
    input [63:0] input_135;
    input [63:0] input_136;
    input [63:0] input_137;
    input [63:0] input_138;
    input [63:0] input_139;
    input [63:0] input_140;
    input [63:0] input_141;
    input [63:0] input_142;
    input [63:0] input_143;
    input [63:0] input_144;
    input [63:0] input_145;
    input [63:0] input_146;
    input [63:0] input_147;
    input [63:0] input_148;
    input [63:0] input_149;
    input [63:0] input_150;
    input [63:0] input_151;
    input [63:0] input_152;
    input [63:0] input_153;
    input [63:0] input_154;
    input [63:0] input_155;
    input [63:0] input_156;
    input [63:0] input_157;
    input [63:0] input_158;
    input [63:0] input_159;
    input [63:0] input_160;
    input [63:0] input_161;
    input [63:0] input_162;
    input [63:0] input_163;
    input [63:0] input_164;
    input [63:0] input_165;
    input [63:0] input_166;
    input [63:0] input_167;
    input [63:0] input_168;
    input [63:0] input_169;
    input [63:0] input_170;
    input [63:0] input_171;
    input [63:0] input_172;
    input [63:0] input_173;
    input [63:0] input_174;
    input [63:0] input_175;
    input [63:0] input_176;
    input [63:0] input_177;
    input [63:0] input_178;
    input [63:0] input_179;
    input [63:0] input_180;
    input [63:0] input_181;
    input [63:0] input_182;
    input [63:0] input_183;
    input [63:0] input_184;
    input [63:0] input_185;
    input [63:0] input_186;
    input [63:0] input_187;
    input [63:0] input_188;
    input [63:0] input_189;
    input [63:0] input_190;
    input [63:0] input_191;
    input [63:0] input_192;
    input [63:0] input_193;
    input [63:0] input_194;
    input [63:0] input_195;
    input [63:0] input_196;
    input [63:0] input_197;
    input [63:0] input_198;
    input [63:0] input_199;
    input [63:0] input_200;
    input [63:0] input_201;
    input [63:0] input_202;
    input [63:0] input_203;
    input [63:0] input_204;
    input [63:0] input_205;
    input [63:0] input_206;
    input [63:0] input_207;
    input [63:0] input_208;
    input [63:0] input_209;
    input [63:0] input_210;
    input [63:0] input_211;
    input [63:0] input_212;
    input [63:0] input_213;
    input [63:0] input_214;
    input [63:0] input_215;
    input [63:0] input_216;
    input [63:0] input_217;
    input [63:0] input_218;
    input [63:0] input_219;
    input [63:0] input_220;
    input [63:0] input_221;
    input [63:0] input_222;
    input [63:0] input_223;
    input [63:0] input_224;
    input [63:0] input_225;
    input [63:0] input_226;
    input [63:0] input_227;
    input [63:0] input_228;
    input [63:0] input_229;
    input [63:0] input_230;
    input [63:0] input_231;
    input [63:0] input_232;
    input [63:0] input_233;
    input [63:0] input_234;
    input [63:0] input_235;
    input [63:0] input_236;
    input [63:0] input_237;
    input [63:0] input_238;
    input [63:0] input_239;
    input [63:0] input_240;
    input [63:0] input_241;
    input [63:0] input_242;
    input [63:0] input_243;
    input [63:0] input_244;
    input [63:0] input_245;
    input [63:0] input_246;
    input [63:0] input_247;
    input [63:0] input_248;
    input [63:0] input_249;
    input [63:0] input_250;
    input [63:0] input_251;
    input [63:0] input_252;
    input [63:0] input_253;
    input [63:0] input_254;
    input [63:0] input_255;
    input [7:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      8'b00000000 : begin
        result = input_0;
      end
      8'b00000001 : begin
        result = input_1;
      end
      8'b00000010 : begin
        result = input_2;
      end
      8'b00000011 : begin
        result = input_3;
      end
      8'b00000100 : begin
        result = input_4;
      end
      8'b00000101 : begin
        result = input_5;
      end
      8'b00000110 : begin
        result = input_6;
      end
      8'b00000111 : begin
        result = input_7;
      end
      8'b00001000 : begin
        result = input_8;
      end
      8'b00001001 : begin
        result = input_9;
      end
      8'b00001010 : begin
        result = input_10;
      end
      8'b00001011 : begin
        result = input_11;
      end
      8'b00001100 : begin
        result = input_12;
      end
      8'b00001101 : begin
        result = input_13;
      end
      8'b00001110 : begin
        result = input_14;
      end
      8'b00001111 : begin
        result = input_15;
      end
      8'b00010000 : begin
        result = input_16;
      end
      8'b00010001 : begin
        result = input_17;
      end
      8'b00010010 : begin
        result = input_18;
      end
      8'b00010011 : begin
        result = input_19;
      end
      8'b00010100 : begin
        result = input_20;
      end
      8'b00010101 : begin
        result = input_21;
      end
      8'b00010110 : begin
        result = input_22;
      end
      8'b00010111 : begin
        result = input_23;
      end
      8'b00011000 : begin
        result = input_24;
      end
      8'b00011001 : begin
        result = input_25;
      end
      8'b00011010 : begin
        result = input_26;
      end
      8'b00011011 : begin
        result = input_27;
      end
      8'b00011100 : begin
        result = input_28;
      end
      8'b00011101 : begin
        result = input_29;
      end
      8'b00011110 : begin
        result = input_30;
      end
      8'b00011111 : begin
        result = input_31;
      end
      8'b00100000 : begin
        result = input_32;
      end
      8'b00100001 : begin
        result = input_33;
      end
      8'b00100010 : begin
        result = input_34;
      end
      8'b00100011 : begin
        result = input_35;
      end
      8'b00100100 : begin
        result = input_36;
      end
      8'b00100101 : begin
        result = input_37;
      end
      8'b00100110 : begin
        result = input_38;
      end
      8'b00100111 : begin
        result = input_39;
      end
      8'b00101000 : begin
        result = input_40;
      end
      8'b00101001 : begin
        result = input_41;
      end
      8'b00101010 : begin
        result = input_42;
      end
      8'b00101011 : begin
        result = input_43;
      end
      8'b00101100 : begin
        result = input_44;
      end
      8'b00101101 : begin
        result = input_45;
      end
      8'b00101110 : begin
        result = input_46;
      end
      8'b00101111 : begin
        result = input_47;
      end
      8'b00110000 : begin
        result = input_48;
      end
      8'b00110001 : begin
        result = input_49;
      end
      8'b00110010 : begin
        result = input_50;
      end
      8'b00110011 : begin
        result = input_51;
      end
      8'b00110100 : begin
        result = input_52;
      end
      8'b00110101 : begin
        result = input_53;
      end
      8'b00110110 : begin
        result = input_54;
      end
      8'b00110111 : begin
        result = input_55;
      end
      8'b00111000 : begin
        result = input_56;
      end
      8'b00111001 : begin
        result = input_57;
      end
      8'b00111010 : begin
        result = input_58;
      end
      8'b00111011 : begin
        result = input_59;
      end
      8'b00111100 : begin
        result = input_60;
      end
      8'b00111101 : begin
        result = input_61;
      end
      8'b00111110 : begin
        result = input_62;
      end
      8'b00111111 : begin
        result = input_63;
      end
      8'b01000000 : begin
        result = input_64;
      end
      8'b01000001 : begin
        result = input_65;
      end
      8'b01000010 : begin
        result = input_66;
      end
      8'b01000011 : begin
        result = input_67;
      end
      8'b01000100 : begin
        result = input_68;
      end
      8'b01000101 : begin
        result = input_69;
      end
      8'b01000110 : begin
        result = input_70;
      end
      8'b01000111 : begin
        result = input_71;
      end
      8'b01001000 : begin
        result = input_72;
      end
      8'b01001001 : begin
        result = input_73;
      end
      8'b01001010 : begin
        result = input_74;
      end
      8'b01001011 : begin
        result = input_75;
      end
      8'b01001100 : begin
        result = input_76;
      end
      8'b01001101 : begin
        result = input_77;
      end
      8'b01001110 : begin
        result = input_78;
      end
      8'b01001111 : begin
        result = input_79;
      end
      8'b01010000 : begin
        result = input_80;
      end
      8'b01010001 : begin
        result = input_81;
      end
      8'b01010010 : begin
        result = input_82;
      end
      8'b01010011 : begin
        result = input_83;
      end
      8'b01010100 : begin
        result = input_84;
      end
      8'b01010101 : begin
        result = input_85;
      end
      8'b01010110 : begin
        result = input_86;
      end
      8'b01010111 : begin
        result = input_87;
      end
      8'b01011000 : begin
        result = input_88;
      end
      8'b01011001 : begin
        result = input_89;
      end
      8'b01011010 : begin
        result = input_90;
      end
      8'b01011011 : begin
        result = input_91;
      end
      8'b01011100 : begin
        result = input_92;
      end
      8'b01011101 : begin
        result = input_93;
      end
      8'b01011110 : begin
        result = input_94;
      end
      8'b01011111 : begin
        result = input_95;
      end
      8'b01100000 : begin
        result = input_96;
      end
      8'b01100001 : begin
        result = input_97;
      end
      8'b01100010 : begin
        result = input_98;
      end
      8'b01100011 : begin
        result = input_99;
      end
      8'b01100100 : begin
        result = input_100;
      end
      8'b01100101 : begin
        result = input_101;
      end
      8'b01100110 : begin
        result = input_102;
      end
      8'b01100111 : begin
        result = input_103;
      end
      8'b01101000 : begin
        result = input_104;
      end
      8'b01101001 : begin
        result = input_105;
      end
      8'b01101010 : begin
        result = input_106;
      end
      8'b01101011 : begin
        result = input_107;
      end
      8'b01101100 : begin
        result = input_108;
      end
      8'b01101101 : begin
        result = input_109;
      end
      8'b01101110 : begin
        result = input_110;
      end
      8'b01101111 : begin
        result = input_111;
      end
      8'b01110000 : begin
        result = input_112;
      end
      8'b01110001 : begin
        result = input_113;
      end
      8'b01110010 : begin
        result = input_114;
      end
      8'b01110011 : begin
        result = input_115;
      end
      8'b01110100 : begin
        result = input_116;
      end
      8'b01110101 : begin
        result = input_117;
      end
      8'b01110110 : begin
        result = input_118;
      end
      8'b01110111 : begin
        result = input_119;
      end
      8'b01111000 : begin
        result = input_120;
      end
      8'b01111001 : begin
        result = input_121;
      end
      8'b01111010 : begin
        result = input_122;
      end
      8'b01111011 : begin
        result = input_123;
      end
      8'b01111100 : begin
        result = input_124;
      end
      8'b01111101 : begin
        result = input_125;
      end
      8'b01111110 : begin
        result = input_126;
      end
      8'b01111111 : begin
        result = input_127;
      end
      8'b10000000 : begin
        result = input_128;
      end
      8'b10000001 : begin
        result = input_129;
      end
      8'b10000010 : begin
        result = input_130;
      end
      8'b10000011 : begin
        result = input_131;
      end
      8'b10000100 : begin
        result = input_132;
      end
      8'b10000101 : begin
        result = input_133;
      end
      8'b10000110 : begin
        result = input_134;
      end
      8'b10000111 : begin
        result = input_135;
      end
      8'b10001000 : begin
        result = input_136;
      end
      8'b10001001 : begin
        result = input_137;
      end
      8'b10001010 : begin
        result = input_138;
      end
      8'b10001011 : begin
        result = input_139;
      end
      8'b10001100 : begin
        result = input_140;
      end
      8'b10001101 : begin
        result = input_141;
      end
      8'b10001110 : begin
        result = input_142;
      end
      8'b10001111 : begin
        result = input_143;
      end
      8'b10010000 : begin
        result = input_144;
      end
      8'b10010001 : begin
        result = input_145;
      end
      8'b10010010 : begin
        result = input_146;
      end
      8'b10010011 : begin
        result = input_147;
      end
      8'b10010100 : begin
        result = input_148;
      end
      8'b10010101 : begin
        result = input_149;
      end
      8'b10010110 : begin
        result = input_150;
      end
      8'b10010111 : begin
        result = input_151;
      end
      8'b10011000 : begin
        result = input_152;
      end
      8'b10011001 : begin
        result = input_153;
      end
      8'b10011010 : begin
        result = input_154;
      end
      8'b10011011 : begin
        result = input_155;
      end
      8'b10011100 : begin
        result = input_156;
      end
      8'b10011101 : begin
        result = input_157;
      end
      8'b10011110 : begin
        result = input_158;
      end
      8'b10011111 : begin
        result = input_159;
      end
      8'b10100000 : begin
        result = input_160;
      end
      8'b10100001 : begin
        result = input_161;
      end
      8'b10100010 : begin
        result = input_162;
      end
      8'b10100011 : begin
        result = input_163;
      end
      8'b10100100 : begin
        result = input_164;
      end
      8'b10100101 : begin
        result = input_165;
      end
      8'b10100110 : begin
        result = input_166;
      end
      8'b10100111 : begin
        result = input_167;
      end
      8'b10101000 : begin
        result = input_168;
      end
      8'b10101001 : begin
        result = input_169;
      end
      8'b10101010 : begin
        result = input_170;
      end
      8'b10101011 : begin
        result = input_171;
      end
      8'b10101100 : begin
        result = input_172;
      end
      8'b10101101 : begin
        result = input_173;
      end
      8'b10101110 : begin
        result = input_174;
      end
      8'b10101111 : begin
        result = input_175;
      end
      8'b10110000 : begin
        result = input_176;
      end
      8'b10110001 : begin
        result = input_177;
      end
      8'b10110010 : begin
        result = input_178;
      end
      8'b10110011 : begin
        result = input_179;
      end
      8'b10110100 : begin
        result = input_180;
      end
      8'b10110101 : begin
        result = input_181;
      end
      8'b10110110 : begin
        result = input_182;
      end
      8'b10110111 : begin
        result = input_183;
      end
      8'b10111000 : begin
        result = input_184;
      end
      8'b10111001 : begin
        result = input_185;
      end
      8'b10111010 : begin
        result = input_186;
      end
      8'b10111011 : begin
        result = input_187;
      end
      8'b10111100 : begin
        result = input_188;
      end
      8'b10111101 : begin
        result = input_189;
      end
      8'b10111110 : begin
        result = input_190;
      end
      8'b10111111 : begin
        result = input_191;
      end
      8'b11000000 : begin
        result = input_192;
      end
      8'b11000001 : begin
        result = input_193;
      end
      8'b11000010 : begin
        result = input_194;
      end
      8'b11000011 : begin
        result = input_195;
      end
      8'b11000100 : begin
        result = input_196;
      end
      8'b11000101 : begin
        result = input_197;
      end
      8'b11000110 : begin
        result = input_198;
      end
      8'b11000111 : begin
        result = input_199;
      end
      8'b11001000 : begin
        result = input_200;
      end
      8'b11001001 : begin
        result = input_201;
      end
      8'b11001010 : begin
        result = input_202;
      end
      8'b11001011 : begin
        result = input_203;
      end
      8'b11001100 : begin
        result = input_204;
      end
      8'b11001101 : begin
        result = input_205;
      end
      8'b11001110 : begin
        result = input_206;
      end
      8'b11001111 : begin
        result = input_207;
      end
      8'b11010000 : begin
        result = input_208;
      end
      8'b11010001 : begin
        result = input_209;
      end
      8'b11010010 : begin
        result = input_210;
      end
      8'b11010011 : begin
        result = input_211;
      end
      8'b11010100 : begin
        result = input_212;
      end
      8'b11010101 : begin
        result = input_213;
      end
      8'b11010110 : begin
        result = input_214;
      end
      8'b11010111 : begin
        result = input_215;
      end
      8'b11011000 : begin
        result = input_216;
      end
      8'b11011001 : begin
        result = input_217;
      end
      8'b11011010 : begin
        result = input_218;
      end
      8'b11011011 : begin
        result = input_219;
      end
      8'b11011100 : begin
        result = input_220;
      end
      8'b11011101 : begin
        result = input_221;
      end
      8'b11011110 : begin
        result = input_222;
      end
      8'b11011111 : begin
        result = input_223;
      end
      8'b11100000 : begin
        result = input_224;
      end
      8'b11100001 : begin
        result = input_225;
      end
      8'b11100010 : begin
        result = input_226;
      end
      8'b11100011 : begin
        result = input_227;
      end
      8'b11100100 : begin
        result = input_228;
      end
      8'b11100101 : begin
        result = input_229;
      end
      8'b11100110 : begin
        result = input_230;
      end
      8'b11100111 : begin
        result = input_231;
      end
      8'b11101000 : begin
        result = input_232;
      end
      8'b11101001 : begin
        result = input_233;
      end
      8'b11101010 : begin
        result = input_234;
      end
      8'b11101011 : begin
        result = input_235;
      end
      8'b11101100 : begin
        result = input_236;
      end
      8'b11101101 : begin
        result = input_237;
      end
      8'b11101110 : begin
        result = input_238;
      end
      8'b11101111 : begin
        result = input_239;
      end
      8'b11110000 : begin
        result = input_240;
      end
      8'b11110001 : begin
        result = input_241;
      end
      8'b11110010 : begin
        result = input_242;
      end
      8'b11110011 : begin
        result = input_243;
      end
      8'b11110100 : begin
        result = input_244;
      end
      8'b11110101 : begin
        result = input_245;
      end
      8'b11110110 : begin
        result = input_246;
      end
      8'b11110111 : begin
        result = input_247;
      end
      8'b11111000 : begin
        result = input_248;
      end
      8'b11111001 : begin
        result = input_249;
      end
      8'b11111010 : begin
        result = input_250;
      end
      8'b11111011 : begin
        result = input_251;
      end
      8'b11111100 : begin
        result = input_252;
      end
      8'b11111101 : begin
        result = input_253;
      end
      8'b11111110 : begin
        result = input_254;
      end
      default : begin
        result = input_255;
      end
    endcase
    MUX_v_64_256_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [15:0] readslicef_27_16_11;
    input [26:0] vector;
    reg [26:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_27_16_11 = tmp[15:0];
  end
  endfunction


  function automatic [10:0] signext_11_1;
    input  vector;
  begin
    signext_11_1= {{10{vector}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input  vector;
  begin
    signext_4_1= {{3{vector}}, vector};
  end
  endfunction


  function automatic [5:0] signext_6_1;
    input  vector;
  begin
    signext_6_1= {{5{vector}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input  vector;
  begin
    signext_7_1= {{6{vector}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [18:0] conv_u2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_u2u_18_19 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore
// ------------------------------------------------------------------


module PECore (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [73:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [96:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [63:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_c;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_en;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_4_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_5_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_6_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_7_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_8_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_9_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_10_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_11_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_12_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_13_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_14_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_15_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_16_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_17_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_18_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_19_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_20_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_b;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_c;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_d;
  wire Datapath_for_4_ProductSum_for_acc_5_cmp_21_en;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_21_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_22_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_23_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_24_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_25_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_26_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_27_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_28_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_29_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_30_z;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_a;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_c;
  wire [17:0] Datapath_for_4_ProductSum_for_acc_5_cmp_31_z;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff;
  wire [7:0] Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_1 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_1_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_1_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_1_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_2 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_2_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_2_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_2_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_3 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_3_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_3_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_3_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_4 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_4_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_4_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_4_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_5 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_5_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_5_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_5_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_6 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_6_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_6_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_6_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_7 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_7_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_7_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_7_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_8 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_8_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_8_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_8_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_9 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_9_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_9_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_9_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_10 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_10_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_10_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_10_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_11 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_11_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_11_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_11_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_12 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_12_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_12_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_12_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_13 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_13_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_13_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_13_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_14 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_14_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_14_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_14_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_15 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_15_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_15_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_15_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_16 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_16_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_16_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_16_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_17 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_17_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_17_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_17_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_18 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_18_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_18_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_18_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_19 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_19_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_19_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_19_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_20 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_20_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_20_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_20_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_21 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_21_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_21_b),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_21_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_21_d),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_21_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_21_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_22 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_22_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_22_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_22_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_23 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_23_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_23_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_23_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_24 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_24_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_24_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_24_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_25 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_25_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_25_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_25_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_26 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_26_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_26_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_26_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_27 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_27_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_27_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_27_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_28 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_28_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_28_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_28_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_29 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_29_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_29_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_29_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_30 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_30_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_30_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_30_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  PECore_mgc_mul2add1_pipe #(.gentype(32'sd1),
  .width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_d(32'sd8),
  .signd_d(32'sd0),
  .width_e(32'sd1),
  .signd_e(32'sd0),
  .width_b2(32'sd0),
  .signd_b2(32'sd0),
  .width_d2(32'sd0),
  .signd_d2(32'sd0),
  .width_z(32'sd18),
  .isadd(32'sd1),
  .add_b2(32'sd1),
  .add_d2(32'sd1),
  .use_const(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd2)) Datapath_for_4_ProductSum_for_acc_5_cmp_31 (
      .a(Datapath_for_4_ProductSum_for_acc_5_cmp_31_a),
      .b(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .c(Datapath_for_4_ProductSum_for_acc_5_cmp_31_c),
      .d(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .cst(1'b0),
      .clk(clk),
      .en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Datapath_for_4_ProductSum_for_acc_5_cmp_31_z),
      .b2(2'b0),
      .d2(2'b0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a0_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a0_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a0_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a0_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a1_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a1_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a1_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_147_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a1_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_PECoreRun PECore_PECoreRun_inst (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_a(Datapath_for_4_ProductSum_for_acc_5_cmp_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_c(Datapath_for_4_ProductSum_for_acc_5_cmp_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_en(Datapath_for_4_ProductSum_for_acc_5_cmp_en),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_z(Datapath_for_4_ProductSum_for_acc_5_cmp_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_a(Datapath_for_4_ProductSum_for_acc_5_cmp_1_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_c(Datapath_for_4_ProductSum_for_acc_5_cmp_1_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_z(Datapath_for_4_ProductSum_for_acc_5_cmp_1_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_a(Datapath_for_4_ProductSum_for_acc_5_cmp_2_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_c(Datapath_for_4_ProductSum_for_acc_5_cmp_2_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_z(Datapath_for_4_ProductSum_for_acc_5_cmp_2_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_a(Datapath_for_4_ProductSum_for_acc_5_cmp_3_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_c(Datapath_for_4_ProductSum_for_acc_5_cmp_3_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_z(Datapath_for_4_ProductSum_for_acc_5_cmp_3_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_4_a(Datapath_for_4_ProductSum_for_acc_5_cmp_4_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_4_c(Datapath_for_4_ProductSum_for_acc_5_cmp_4_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_4_z(Datapath_for_4_ProductSum_for_acc_5_cmp_4_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_a(Datapath_for_4_ProductSum_for_acc_5_cmp_5_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_c(Datapath_for_4_ProductSum_for_acc_5_cmp_5_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_5_z(Datapath_for_4_ProductSum_for_acc_5_cmp_5_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_6_a(Datapath_for_4_ProductSum_for_acc_5_cmp_6_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_6_c(Datapath_for_4_ProductSum_for_acc_5_cmp_6_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_6_z(Datapath_for_4_ProductSum_for_acc_5_cmp_6_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_7_a(Datapath_for_4_ProductSum_for_acc_5_cmp_7_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_7_c(Datapath_for_4_ProductSum_for_acc_5_cmp_7_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_7_z(Datapath_for_4_ProductSum_for_acc_5_cmp_7_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_8_a(Datapath_for_4_ProductSum_for_acc_5_cmp_8_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_8_c(Datapath_for_4_ProductSum_for_acc_5_cmp_8_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_8_z(Datapath_for_4_ProductSum_for_acc_5_cmp_8_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_9_a(Datapath_for_4_ProductSum_for_acc_5_cmp_9_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_9_c(Datapath_for_4_ProductSum_for_acc_5_cmp_9_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_9_z(Datapath_for_4_ProductSum_for_acc_5_cmp_9_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_10_a(Datapath_for_4_ProductSum_for_acc_5_cmp_10_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_10_c(Datapath_for_4_ProductSum_for_acc_5_cmp_10_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_10_z(Datapath_for_4_ProductSum_for_acc_5_cmp_10_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_11_a(Datapath_for_4_ProductSum_for_acc_5_cmp_11_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_11_c(Datapath_for_4_ProductSum_for_acc_5_cmp_11_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_11_z(Datapath_for_4_ProductSum_for_acc_5_cmp_11_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_12_a(Datapath_for_4_ProductSum_for_acc_5_cmp_12_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_12_c(Datapath_for_4_ProductSum_for_acc_5_cmp_12_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_12_z(Datapath_for_4_ProductSum_for_acc_5_cmp_12_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_13_a(Datapath_for_4_ProductSum_for_acc_5_cmp_13_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_13_c(Datapath_for_4_ProductSum_for_acc_5_cmp_13_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_13_z(Datapath_for_4_ProductSum_for_acc_5_cmp_13_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_14_a(Datapath_for_4_ProductSum_for_acc_5_cmp_14_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_14_c(Datapath_for_4_ProductSum_for_acc_5_cmp_14_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_14_z(Datapath_for_4_ProductSum_for_acc_5_cmp_14_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_15_a(Datapath_for_4_ProductSum_for_acc_5_cmp_15_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_15_c(Datapath_for_4_ProductSum_for_acc_5_cmp_15_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_15_z(Datapath_for_4_ProductSum_for_acc_5_cmp_15_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_16_a(Datapath_for_4_ProductSum_for_acc_5_cmp_16_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_16_c(Datapath_for_4_ProductSum_for_acc_5_cmp_16_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_16_z(Datapath_for_4_ProductSum_for_acc_5_cmp_16_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_17_a(Datapath_for_4_ProductSum_for_acc_5_cmp_17_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_17_c(Datapath_for_4_ProductSum_for_acc_5_cmp_17_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_17_z(Datapath_for_4_ProductSum_for_acc_5_cmp_17_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_18_a(Datapath_for_4_ProductSum_for_acc_5_cmp_18_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_18_c(Datapath_for_4_ProductSum_for_acc_5_cmp_18_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_18_z(Datapath_for_4_ProductSum_for_acc_5_cmp_18_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_19_a(Datapath_for_4_ProductSum_for_acc_5_cmp_19_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_19_c(Datapath_for_4_ProductSum_for_acc_5_cmp_19_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_19_z(Datapath_for_4_ProductSum_for_acc_5_cmp_19_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_20_a(Datapath_for_4_ProductSum_for_acc_5_cmp_20_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_20_c(Datapath_for_4_ProductSum_for_acc_5_cmp_20_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_20_z(Datapath_for_4_ProductSum_for_acc_5_cmp_20_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_a(Datapath_for_4_ProductSum_for_acc_5_cmp_21_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_b(Datapath_for_4_ProductSum_for_acc_5_cmp_21_b),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_c(Datapath_for_4_ProductSum_for_acc_5_cmp_21_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_d(Datapath_for_4_ProductSum_for_acc_5_cmp_21_d),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_en(Datapath_for_4_ProductSum_for_acc_5_cmp_21_en),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_21_z(Datapath_for_4_ProductSum_for_acc_5_cmp_21_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_22_a(Datapath_for_4_ProductSum_for_acc_5_cmp_22_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_22_c(Datapath_for_4_ProductSum_for_acc_5_cmp_22_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_22_z(Datapath_for_4_ProductSum_for_acc_5_cmp_22_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_23_a(Datapath_for_4_ProductSum_for_acc_5_cmp_23_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_23_c(Datapath_for_4_ProductSum_for_acc_5_cmp_23_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_23_z(Datapath_for_4_ProductSum_for_acc_5_cmp_23_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_24_a(Datapath_for_4_ProductSum_for_acc_5_cmp_24_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_24_c(Datapath_for_4_ProductSum_for_acc_5_cmp_24_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_24_z(Datapath_for_4_ProductSum_for_acc_5_cmp_24_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_25_a(Datapath_for_4_ProductSum_for_acc_5_cmp_25_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_25_c(Datapath_for_4_ProductSum_for_acc_5_cmp_25_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_25_z(Datapath_for_4_ProductSum_for_acc_5_cmp_25_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_26_a(Datapath_for_4_ProductSum_for_acc_5_cmp_26_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_26_c(Datapath_for_4_ProductSum_for_acc_5_cmp_26_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_26_z(Datapath_for_4_ProductSum_for_acc_5_cmp_26_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_27_a(Datapath_for_4_ProductSum_for_acc_5_cmp_27_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_27_c(Datapath_for_4_ProductSum_for_acc_5_cmp_27_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_27_z(Datapath_for_4_ProductSum_for_acc_5_cmp_27_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_28_a(Datapath_for_4_ProductSum_for_acc_5_cmp_28_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_28_c(Datapath_for_4_ProductSum_for_acc_5_cmp_28_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_28_z(Datapath_for_4_ProductSum_for_acc_5_cmp_28_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_29_a(Datapath_for_4_ProductSum_for_acc_5_cmp_29_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_29_c(Datapath_for_4_ProductSum_for_acc_5_cmp_29_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_29_z(Datapath_for_4_ProductSum_for_acc_5_cmp_29_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_30_a(Datapath_for_4_ProductSum_for_acc_5_cmp_30_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_30_c(Datapath_for_4_ProductSum_for_acc_5_cmp_30_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_30_z(Datapath_for_4_ProductSum_for_acc_5_cmp_30_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_31_a(Datapath_for_4_ProductSum_for_acc_5_cmp_31_a),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_31_c(Datapath_for_4_ProductSum_for_acc_5_cmp_31_c),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_31_z(Datapath_for_4_ProductSum_for_acc_5_cmp_31_z),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_1_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_1_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_2_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_2_d_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_3_b_iff),
      .Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_pff(Datapath_for_4_ProductSum_for_acc_5_cmp_3_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff)
    );
endmodule



